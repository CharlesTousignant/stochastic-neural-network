library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;
use ieee.numeric_std.all;
use IEEE.math_real.all; 

package utilsAxiWrapper is
    type pixelVec is array(783 downto 0) of unsigned(33 downto 0);
end package;

package body utilsAxiWrapper is
  
end package body;