library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;  	
use work.all;
use work.utils.all;

entity LFSR is 
    generic(seed: integer);
    port (
	clk, reset : in std_logic;
    random: out std_logic_vector(31 downto 0)
	);
end LFSR;
-- esrer dwdawdw
architecture arch of LFSR is	
constant seed1: std_logic_vector(63 downto 0) := std_logic_vector(rand_slv(64, (seed - 1) * 3 + 1));
constant differentTaps: LFSRPolynomial := 
(x"800000000000000D",
 x"800000000000000E",
 x"800000000000007A",
 x"80000000000000BA",
 x"80000000000000D0",
 x"80000000000000EF",
 x"8000000000000128",
 x"8000000000000165",
 x"80000000000001A3",
 x"80000000000001E4",
 x"80000000000001E7",
 x"80000000000001F9",
 x"8000000000000212",
 x"8000000000000299",
 x"80000000000003BC",
 x"80000000000003BF",
 x"8000000000000403",
 x"8000000000000472",
 x"800000000000049C",
 x"80000000000004C9",
 x"8000000000000508",
 x"800000000000056B",
 x"800000000000057C",
 x"8000000000000645",
 x"8000000000000658",
 x"8000000000000703",
 x"8000000000000711",
 x"8000000000000784",
 x"80000000000007B4",
 x"80000000000007C9",
 x"80000000000007F5",
 x"8000000000000841",
 x"8000000000000869",
 x"800000000000089C",
 x"80000000000008F6",
 x"8000000000000940",
 x"8000000000000952",
 x"8000000000000957",
 x"800000000000096D",
 x"8000000000000B22",
 x"8000000000000B24",
 x"8000000000000B2D",
 x"8000000000000B44",
 x"8000000000000B84",
 x"8000000000000BA3",
 x"8000000000000BAF",
 x"8000000000000BC3",
 x"8000000000000CBC",
 x"8000000000000D0F",
 x"8000000000000D18",
 x"8000000000000D27",
 x"8000000000000D71",
 x"8000000000000DAA",
 x"8000000000000DDD",
 x"8000000000000E2E",
 x"8000000000000E5C",
 x"8000000000000E82",
 x"8000000000000EB7",
 x"8000000000000EC3",
 x"8000000000000EFA",
 x"8000000000000FC1",
 x"8000000000000FE3",
 x"800000000000101B",
 x"800000000000102B",
 x"8000000000001036",
 x"80000000000010CA",
 x"80000000000010F0",
 x"800000000000114C",
 x"800000000000115E",
 x"800000000000117F",
 x"80000000000011D5",
 x"80000000000011E5",
 x"8000000000001237",
 x"8000000000001238",
 x"800000000000125E",
 x"80000000000012DF",
 x"8000000000001324",
 x"8000000000001335",
 x"8000000000001395",
 x"8000000000001410",
 x"800000000000143D",
 x"800000000000147C",
 x"80000000000014C1",
 x"80000000000014F8",
 x"800000000000155C",
 x"80000000000015B7",
 x"80000000000015D1",
 x"8000000000001618",
 x"8000000000001713",
 x"8000000000001797",
 x"80000000000017AE",
 x"8000000000001858",
 x"8000000000001868",
 x"80000000000018F8",
 x"8000000000001933",
 x"800000000000193A",
 x"800000000000196C",
 x"800000000000198B",
 x"80000000000019A9",
 x"80000000000019E2"
);
constant chosenTaps : std_logic_vector (63 downto 0) :=  differentTaps( to_integer(unsigned(seed1) mod 100));
signal state : std_logic_vector (63 downto 0) :=  seed1;
begin	
						    
    process(clk)
    variable newBit: std_logic;
    begin
    if (rising_edge(clk)) then
    
        if(reset = '1') then
            state <= seed1;
        else    
            newBit := xor(state and chosenTaps);
            state <= state(62 downto 0) & newBit;
        end if;
    end if;
	end process;
	
	random <= state(63 downto 32);
end arch;