library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;
use ieee.numeric_std.all;
use IEEE.math_real.all; 

package utils is
    constant precision: integer := 10; -- the precision in number of bits, stream length = 2**precision
    constant m : integer := 1;
    -- constant mPrime : integer := 6;
    
    type neuronWeights is array(natural range <>) of std_logic_vector(31 downto 0);
    subtype neuronBias is std_logic_vector(31 downto 0);
	
	type randomNumberVector is array(natural range <>) of std_logic_vector(31 downto 0);
    type layerWeights is array(natural range <>) of neuronWeights; 
    type layerBiases is array(natural range <>) of neuronBias;
    type layerScales is array(natural range<>) of integer;
    
    type networkInputs is array(natural range<>) of std_logic_vector (31 downto 0);  
    type networkInputsArray10 is array(natural range<>) of networkInputs(0 to 9);
    type networkInputsArray is array(natural range<>) of networkInputs(0 to 783);
    type networkExpectedOuputs is array(natural range<>) of natural;
    
    subtype neuronOutput is std_logic_vector (precision - 1 downto 0);
    type networkOutputs is array(natural range <>) of neuronOutput;
    
    type LFSRPolynomial is array(natural range<>) of std_logic_vector;
	
    function f_log2 (x: positive) return natural;
    function muxSelectFromRand(rand: std_logic_vector(31 downto 0); numEntries: integer) return integer;
	function bitAdderTree(v: std_logic_vector) return natural;

    type CTStateValue is array(2 downto 0) of unsigned(31 downto 0);
    type CTState is protected
      -- Definition of functions and procedures
      procedure set(newState: CTStateValue);
      impure function get_value return CTStateValue;
    end protected CTState;

    impure function rand_slv(len : integer; seed : integer) return unsigned;
    type randSeeds is array(7065 downto 1) of std_logic_vector(31 downto 0);
    constant seeds: randSeeds := (x"d091bb5c" , x"22ae9ef6" , x"e7e1faee" , x"d5c31f79" , x"2082352c" , x"f807b7df" , x"e9d30005" , x"3895afe1" , x"a1e24bba" , x"4ee4092b" , x"18f86863" , x"8c16a625" , x"474ba8c4" , x"3039cd1a" , x"8c006d5f" , x"fe2d7810" , x"f51f2ae7" , x"ff1816e4" , x"f702ef59" , x"f7badafa" , x"285954a1" , x"b9d09511" , x"f878c4b3" , x"fb2a0137" , x"f508e4aa" , x"1c1fe652" , x"7c419418" , x"cc50aa59" , x"ccdf2e5c" , x"4c0a1f3b" , x"2452a9dc" , x"01397d8d" , x"6bf88c31" , x"1cca797a" , x"ea6da4ae" , x"a3c78807" , x"cace1969" , x"e0e0d4ad" , x"f5a14bab" , x"80f00988" , x"a7de9f4c" , x"cc450cba" , x"0924668f" , x"5c7dc380" , x"d96089c5" , x"3640ac4c" , x"ef1a2e6d" , x"ae6d9426" , x"adc1965b" , x"6613ba46" , x"c1fb41c2" , x"bd9b0ecd" , x"be3dedfc" , x"7989c8ee" , x"6468fd6e" , x"6c0df032" , x"a7cd6634" , x"2c826d8b" , x"2bd2e412" , x"4d4a2dbe" , x"b4bf6fa7" , x"cc1a8959" , x"08263282" , x"51097330" , x"46e46cb0" , x"df577ec2" , x"0bd1e364" , x"262c5564" , x"18dda0c9" , x"fe7b45d9" , x"d2ce21c9" , x"d268409a" , x"b1e049e1" , x"200bfa47" , x"512d6e73" , x"c3851eee" , x"f341c081" , x"7d973e48" , x"08d17554" , x"a9e20d28" , x"70518ce6" , x"203ac303" , x"61add0ab" , x"35d0430c" , x"c3f8e892" , x"0d1c8509" , x"cb92388e" , x"095436bf" , x"2fd6e208" , x"68a29af9" , x"7d61330b" , x"753ec6fc" , x"7211efea" , x"7cd15133" , x"a574c4ff" , x"cb41f198" , x"b598eef6" , x"ebbe7347" , x"c1332568" , x"ceba5a70" , x"46a99459" , x"b4ad9f11" , x"ae00feaa" , x"00b8b573" , x"a7b480b6" , x"b5f0b06c" , x"29a0ec27" , x"a4daa010" , x"1e76a1c5" , x"74be9133" , x"7f94c950" , x"c61f6ed6" , x"f5b1c7a1" , x"92e195f8" , x"572384d4" , x"e0732c88" , x"95d41b68" , x"cee496c3" , x"394bbd52" , x"048cd47c" , x"c05309be" , x"d23d2d63" , x"414de9c5" , x"d2229f23" , x"818666a3" , x"f0a8b109" , x"b2f6b127" , x"69a48341" , x"e4123c56" , x"6c548c8f" , x"f5941f61" , x"94b993aa" , x"8c165134" , x"2876763c" , x"237ce42e" , x"c300d11b" , x"263821ca" , x"3aeb8202" , x"41ec0f84" , x"cf4ac36d" , x"d7393ee6" , x"fd0fc06a" , x"4118a30a" , x"551b54a4" , x"d074f86f" , x"4cc1c54a" , x"3e57a703" , x"03774cda" , x"ede43895" , x"379ce627" , x"59988939" , x"e8490ddc" , x"325410e1" , x"d9352f6a" , x"4047080a" , x"f47c081d" , x"9db51a85" , x"c765d71f" , x"79297527" , x"fcca2773" , x"5a065b97" , x"114dee4f" , x"d4b12f5f" , x"cb29360a" , x"95d3de16" , x"983162a8" , x"8cbaafb3" , x"bb98b27f" , x"eacd3439" , x"b1fac842" , x"492cbef1" , x"ae08ab78" , x"c1d7dfd0" , x"646f1d40" , x"c0f463c4" , x"8fc23a81" , x"6164e623" , x"3543f2bc" , x"915cc253" , x"8701d0df" , x"136b2fdd" , x"677a359e" , x"0dcfacd0" , x"5a4ea31e" , x"87e25935" , x"97c34e42" , x"c77780f0" , x"5b396fba" , x"ef1b52e6" , x"f7080941" , x"2141888b" , x"278946b0" , x"919e6d64" , x"6518b459" , x"7829fc22" , x"6325d30e" , x"030c0399" , x"ba19b463" , x"564dab75" , x"63794f97" , x"2984c787" , x"ed702bbe" , x"cb563b4d" , x"6fa56696" , x"4fabc9ed" , x"dcd87a48" , x"874df295" , x"9ecfe9f0" , x"2a67f49f" , x"1e9aa4e1" , x"9a1b7d08" , x"78d22934" , x"43521602" , x"5718a361" , x"a771ba44" , x"87a3b97c" , x"b0705c82" , x"b7526048" , x"bf86dcd7" , x"fd066ea4" , x"7356b1bb" , x"b872426d" , x"1575515d" , x"e99eadb3" , x"3a9e3c0f" , x"8168599c" , x"e9d07a32" , x"8eeab382" , x"27023ee8" , x"80d10fac" , x"d368bdc2" , x"7664b5a7" , x"89d0cf46" , x"8bed7368" , x"ff02af49" , x"7294e430" , x"14034fbb" , x"dabd4cc4" , x"71535cf8" , x"9aaeea20" , x"1b4d989d" , x"7fa09780" , x"f63ef3d2" , x"fadc6788" , x"012fb568" , x"08c904fa" , x"c660883f" , x"fa1cce2a" , x"d13ac8b8" , x"5cf9c9b3" , x"de62c6bd" , x"adf500ad" , x"159d967e" , x"58a2c06c" , x"665827cb" , x"db1aa208" , x"4286ddf1" , x"0b8905b4" , x"ccd149a4" , x"a8fd9757" , x"6e7122f0" , x"bffc21b1" , x"e9203368" , x"220c0724" , x"2e8d86cb" , x"fb7bfb5e" , x"43889687" , x"1869325b" , x"25420afc" , x"485d46db" , x"22d56381" , x"cd572d60" , x"de89ef2b" , x"13dac708" , x"9467851d" , x"a09c428d" , x"8cc3a36c" , x"0212714e" , x"251bc1f6" , x"ae274af0" , x"da603f48" , x"88afd714" , x"9f3f014d" , x"704c7830" , x"59d803fb" , x"3315c9dc" , x"83645273" , x"23540e0e" , x"66dce437" , x"61e09244" , x"13728d90" , x"c32e0a94" , x"3d6b2529" , x"0a5c5094" , x"1f91d464" , x"40c1b904" , x"2f1494b9" , x"8138ac02" , x"3d6d8755" , x"d2963cf5" , x"6ad203b6" , x"fb5234e0" , x"0cb62703" , x"d2cdf95b" , x"e718672d" , x"4d448df1" , x"f1dd92d7" , x"0c4613a1" , x"7da944f1" , x"3f72f0c3" , x"7d3fa930" , x"8b4742bc" , x"5674c771" , x"e3420514" , x"e669edd5" , x"5805de29" , x"5e86f504" , x"088449f4" , x"1c77c8a0" , x"29b1fccc" , x"c7be9961" , x"e09aebe7" , x"63c5ecb9" , x"35d657e1" , x"3ddf7ae4" , x"45d3249c" , x"6766c940" , x"7e10ad9c" , x"18b13e7f" , x"39320ca2" , x"21c90078" , x"7d84661c" , x"f12a3a21" , x"f4772b41" , x"f4c53bab" , x"a6e76b3b" , x"9340ded2" , x"c1ebc21f" , x"0f4db654" , x"6f6c42e3" , x"3c1a8943" , x"8d899f74" , x"5a6899ba" , x"0d9b6827" , x"d239c5cb" , x"5290106a" , x"03f17adb" , x"67acdc26" , x"0b039b90" , x"e88f1afa" , x"2b42ee31" , x"cf239e4d" , x"a62c6e93" , x"421fae11" , x"bb522891" , x"213d9f32" , x"a5d2adeb" , x"7e4aab21" , x"736fbc75" , x"60e56773" , x"8c08c64d" , x"b7eda589" , x"4bdbae33" , x"49ad9663" , x"bea4300c" , x"9f997956" , x"305f5b0c" , x"cfd6f924" , x"afd083db" , x"500085e0" , x"2efa9644" , x"62bdecbd" , x"5e5501a5" , x"580bc7bb" , x"a02889ad" , x"d0d63dcd" , x"c7bcfc3c" , x"ab56454f" , x"14c4a882" , x"612197c7" , x"edec3d2f" , x"75600d88" , x"c6951b28" , x"4db9a52d" , x"7c9e604d" , x"e91ac974" , x"6f946da2" , x"7d160cf0" , x"72606b78" , x"c17b7257" , x"4e6ceb4e" , x"1ba9f219" , x"822d9f9a" , x"64c24df6" , x"82c1eccb" , x"dec48f52" , x"d1500cb6" , x"5c615e22" , x"cb7a1247" , x"eac83d5e" , x"a4f2087e" , x"8b36d663" , x"60ec8b7d" , x"23e07770" , x"cfc3bcb6" , x"332ade50" , x"886741fc" , x"f2ecc125" , x"59c94057" , x"fd77d893" , x"f062680f" , x"3d759e10" , x"e03dc9c3" , x"043ab169" , x"8cd70bce" , x"637c48af" , x"9f5a86f9" , x"c799b8ed" , x"96488fc2" , x"7a04f3e1" , x"352e9955" , x"8a467bfe" , x"4d1e7adb" , x"04b931c9" , x"788e6ea0" , x"e67267f5" , x"3b0145b6" , x"31ca7310" , x"d8249eec" , x"e2d0c5d1" , x"31dc1298" , x"70f4055d" , x"39d60297" , x"25d81f3b" , x"2bb385c9" , x"3d500890" , x"3a48350d" , x"ccb6120b" , x"6f89f2f9" , x"791783d6" , x"4fa4664e" , x"16fea67f" , x"ec629bbf" , x"a5014386" , x"6e221244" , x"a21075d9" , x"2f501f52" , x"959a12f4" , x"e7a64774" , x"ba060582" , x"fad0ca2f" , x"5ac9908f" , x"7059c853" , x"ae2f213e" , x"1c724f28" , x"b51305fc" , x"42108734" , x"298e5c9d" , x"68a1dd2b" , x"223c8c36" , x"984b1bef" , x"73161b54" , x"43204f20" , x"0ac40f25" , x"9a53eca9" , x"cc200dd8" , x"b6123cc0" , x"2ae4efad" , x"38c464c2" , x"d4ca75a4" , x"1e0f1559" , x"5330cf6e" , x"4bf2f32b" , x"a7e130fd" , x"519b7462" , x"6b919194" , x"6c963148" , x"c82b32bb" , x"82030024" , x"1cfa2fa0" , x"15e45ce2" , x"fe584a91" , x"4332093f" , x"2e7b9117" , x"cd0f4b4d" , x"c34f792c" , x"077afaf5" , x"44136041" , x"edc96297" , x"3e7fd864" , x"baf6f6ba" , x"19c9ff6e" , x"7d157a58" , x"5825dfde" , x"941a37e0" , x"4818babb" , x"3cbe9dc1" , x"f7f8d0ce" , x"75771de9" , x"36b9cf69" , x"f68cf878" , x"9b1e1c75" , x"8bfb75ae" , x"39ff446d" , x"85692875" , x"309da59f" , x"3b49c509" , x"66cd636e" , x"7d286708" , x"69cd6a2e" , x"9fc266e3" , x"2b8f1988" , x"addbd3af" , x"4c8ea8e7" , x"65407c37" , x"a2ef9aa6" , x"5e10541b" , x"26cd9065" , x"fcec6367" , x"c4ed1ef8" , x"09a9410f" , x"e24bc427" , x"e29a5edd" , x"f58f8c10" , x"e9cd2a63" , x"049ffdb7" , x"cbd2b4cc" , x"95356bb0" , x"19453535" , x"c4508ca2" , x"4309fd7e" , x"53ea8de9" , x"55d9f238" , x"210a7aea" , x"ae02a6ab" , x"4abdf123" , x"22f5256b" , x"d8dc2d8e" , x"b8a25d9d" , x"3b13600f" , x"1b54beda" , x"808164b1" , x"a75ca457" , x"0068b861" , x"7e822ee1" , x"0335be36" , x"c76fef0e" , x"495dbce8" , x"b70cab9d" , x"19445725" , x"e75a3b16" , x"627f5136" , x"e4137f41" , x"5af821c1" , x"558bb5a6" , x"b85003e7" , x"b2e101c2" , x"10c101fc" , x"32a3aa3d" , x"838c4690" , x"07d18800" , x"6c89d813" , x"be7ba68d" , x"b096d0b9" , x"8001786a" , x"41026a58" , x"7adc2d65" , x"66c9fc5f" , x"e79be068" , x"43b4bc3b" , x"9c203868" , x"ef2b0be2" , x"9e1f6267" , x"78f76a0a" , x"dc04692d" , x"9c6500f3" , x"ce348e12" , x"7d07e7ee" , x"93a40579" , x"83b78de9" , x"2ed401c8" , x"3eb994dd" , x"3d6c2f3d" , x"553fd4da" , x"e2f27231" , x"809ad218" , x"0757306e" , x"989740b3" , x"7d6a2d71" , x"4f66622b" , x"2afd45f7" , x"f687016b" , x"fa8ad0b3" , x"3b7e96f2" , x"b6732508" , x"bf351d33" , x"801ee898" , x"5291851f" , x"78993f7e" , x"5177a95e" , x"0f432e84" , x"f3d5350c" , x"ae95b5e0" , x"88e37a7b" , x"0adcc451" , x"df2e9f5b" , x"124a3fe8" , x"ef421e88" , x"858ad803" , x"aac7fd11" , x"18c34c95" , x"4a2915bb" , x"d1722f1a" , x"10c6360b" , x"d14ac42f" , x"3b5d0d66" , x"b8f1cd0d" , x"b468c613" , x"265d94fd" , x"31f28f03" , x"a8dbe3dd" , x"6c16811b" , x"84c2a353" , x"efa14dff" , x"f914dc58" , x"246858c1" , x"a6244e68" , x"a4a782a4" , x"cce276f9" , x"7904f936" , x"742c1628" , x"6fdad5d1" , x"6eb135b6" , x"3e8bbb60" , x"d347c3df" , x"8183ef4e" , x"155e4713" , x"e82d7cf3" , x"22177ec5" , x"1395c3b0" , x"2c633227" , x"b6c26847" , x"64147fff" , x"9e012434" , x"d4d54d85" , x"3067d25f" , x"cda949fd" , x"65a09982" , x"0f7b0a12" , x"4714fddd" , x"6635c1c5" , x"dbac6554" , x"86e1558d" , x"e8b0113e" , x"6ab35ea6" , x"9e06008a" , x"a827f848" , x"2e4a226e" , x"a0c2dcab" , x"83d89830" , x"4abf77e8" , x"d31b1042" , x"6e80b0f7" , x"5bfcafb4" , x"03f6f6ce" , x"d0ed0b8a" , x"fbeb99af" , x"4b1b7def" , x"2acb8c9c" , x"2c0fe9b1" , x"1b30fe94" , x"7e277559" , x"5f563ea0" , x"3200cdd8" , x"32b7e32a" , x"dd43417d" , x"7d5c2b5b" , x"344643f9" , x"56e90a5f" , x"9dc40517" , x"f39e0dc7" , x"e0c7ebbf" , x"eb9ae161" , x"6478daa3" , x"0d7c3d4e" , x"f252e312" , x"bce444b9" , x"2aacbcdb" , x"44e502aa" , x"f8ccf513" , x"6c3ef465" , x"906000da" , x"8c41446a" , x"992eb47b" , x"f1573608" , x"2197c153" , x"6af14701" , x"911852c9" , x"fba9538f" , x"8debdd8c" , x"4d2c26d1" , x"4f7c4522" , x"b37b354f" , x"1ee2d92c" , x"aa952ed2" , x"bcdfdbf3" , x"8a043123" , x"3e232325" , x"b2b70b0d" , x"d2a6e5a6" , x"aaa192d4" , x"2f7b5a6e" , x"2d9a16b1" , x"500b9889" , x"20c58d24" , x"e1b8c1bc" , x"ffc3bb81" , x"ac993839" , x"2bce9702" , x"bd429acc" , x"08588715" , x"1002d574" , x"8faaca38" , x"21ae04bc" , x"e1c200dd" , x"17072760" , x"ab4f12b3" , x"0220e53e" , x"30c03c0a" , x"74ddddc9" , x"5e71509d" , x"a261b3d2" , x"75f22283" , x"879e8c26" , x"fb4c9fe6" , x"7f745ef0" , x"280a27b6" , x"55f6d9e0" , x"db038ae1" , x"40b907f0" , x"a50f49f3" , x"3bd2275a" , x"6053602f" , x"2c546996" , x"30e06018" , x"9892367a" , x"6da1fcf7" , x"ba15ab48" , x"7b65cc3d" , x"e0a8a155" , x"1ee06716" , x"b5086b7b" , x"96e9f667" , x"3c19993c" , x"39e76f8f" , x"7a5dede2" , x"62766632" , x"04a986ae" , x"953e9871" , x"bf5118f1" , x"40765da0" , x"a79bf6f2" , x"4a5a51cc" , x"13fc31f4" , x"9df9ab13" , x"79076552" , x"43e97309" , x"ff18fd70" , x"d30a52a7" , x"88378b0f" , x"fb8fd412" , x"e6417027" , x"baf195a7" , x"c5dcd5cd" , x"580852da" , x"3429986e" , x"95859146" , x"e838454a" , x"1b96c004" , x"5ff3b74d" , x"e803cf9c" , x"d91c5a75" , x"e130fc96" , x"53a28fd0" , x"d158c194" , x"53a50385" , x"42bf11f5" , x"a8c206f5" , x"9827bb23" , x"96363ad9" , x"05c362a9" , x"0c8a29c4" , x"6cddcb78" , x"c51c7848" , x"500e585a" , x"7de37864" , x"2957106e" , x"7cf9a0ab" , x"2dc39ee9" , x"6ddb3d2b" , x"6c423c98" , x"650ce024" , x"181f69eb" , x"c6c5ad24" , x"9938d8c1" , x"f98980e3" , x"788e7de8" , x"bf9e08bc" , x"b229bbe9" , x"a26eb92b" , x"b32bd9ac" , x"127a67ca" , x"a376c062" , x"a22418d6" , x"089a42d0" , x"876757b3" , x"119d46da" , x"4bd1a4a8" , x"51d149d4" , x"5348afee" , x"87e6b8af" , x"a191134a" , x"a789c0f8" , x"fe97e849" , x"6859bb5c" , x"841bb5db" , x"d1ea4a06" , x"b975cfca" , x"b7e65f3f" , x"3eddfc98" , x"f7f96715" , x"55142d20" , x"88057fbb" , x"bfa4d8d4" , x"533cbf5e" , x"aed6e43f" , x"1b0a83f1" , x"ae67ccf0" , x"9c67c962" , x"142f0382" , x"c75f956a" , x"757cd939" , x"6c67691a" , x"b2b9c0a8" , x"174031e8" , x"1160e67b" , x"443779d1" , x"11b3299a" , x"27560be1" , x"86ec4732" , x"47eff6b9" , x"4315a14c" , x"70a96b74" , x"7bbe7982" , x"86f2d3ae" , x"217c7787" , x"7519c371" , x"182d452c" , x"e0185a62" , x"1ed1557a" , x"849f1010" , x"f8474049" , x"f1914086" , x"c19bac85" , x"a340e755" , x"44a73507" , x"f52b6e09" , x"b9937043" , x"3d9ef9f4" , x"6a6f6972" , x"ad1659e7" , x"7987252a" , x"4a0022c0" , x"0e3168c9" , x"abfb9eb5" , x"9d1e560e" , x"b1f4ba47" , x"7d993809" , x"1167f948" , x"e78baa36" , x"4139ed77" , x"ef6a33d1" , x"395aafe9" , x"eb142d32" , x"aaf715e6" , x"4dc77e33" , x"d82a1596" , x"ca441c2b" , x"582eb04f" , x"39ea0a16" , x"c7d022df" , x"72ee825e" , x"ace28fef" , x"82967f6a" , x"01b81854" , x"3b0ab1a1" , x"9a27d844" , x"b63dd19c" , x"63036fc5" , x"fc051613" , x"ea7e66eb" , x"a7bc0e30" , x"004b6f8a" , x"45cd80de" , x"76631166" , x"78116769" , x"6ca2239f" , x"00c4afde" , x"75fe9d74" , x"7248d6c0" , x"c5293013" , x"f88fcbbb" , x"528d833b" , x"4dfe6d59" , x"c8e4aca6" , x"371162e7" , x"78aadccb" , x"3f61bc3b" , x"0927bf11" , x"ce739311" , x"2d061b1e" , x"7c82d0fa" , x"b8c52266" , x"68520ba8" , x"793660d8" , x"37337b3e" , x"2718bc8d" , x"8a4df5f5" , x"5753f130" , x"b9181dce" , x"9b7ddc13" , x"48a02a1b" , x"31163787" , x"8af902aa" , x"bd098a99" , x"c18447b7" , x"3e2b642e" , x"54fc76a4" , x"eadc525a" , x"cd405695" , x"44e13850" , x"db691951" , x"c3f7cf36" , x"03cff145" , x"304c26ac" , x"e28b9a3e" , x"49997af9" , x"97d48bb6" , x"17533654" , x"16125513" , x"9382753b" , x"ecc4ab75" , x"aef0e4a3" , x"e9e9869f" , x"8bed86b3" , x"fb12e042" , x"6cfc90a6" , x"e667d955" , x"a4fa33b5" , x"f3207eb6" , x"a5ca44c1" , x"ef3cd4b0" , x"add40ac4" , x"02218a17" , x"a2c2eaef" , x"c71d8276" , x"f1f6ee43" , x"06a53db2" , x"357cc25f" , x"967f1c3e" , x"b5937c41" , x"a6580857" , x"3c799b6c" , x"54074de7" , x"1e90c0a2" , x"1c6fb273" , x"9b78456a" , x"1fd05538" , x"733c3941" , x"f9527f4f" , x"756f08b1" , x"8881ba01" , x"a975360d" , x"a98c82e2" , x"c5316e71" , x"b5505f48" , x"59a7e348" , x"1198da00" , x"a9797612" , x"34b98139" , x"6a895e81" , x"6ef53f4e" , x"d788ab48" , x"02dd8470" , x"d53a0971" , x"11bb305a" , x"41a61df7" , x"57d2e616" , x"9d0bc340" , x"4fee4f80" , x"950e47fd" , x"fe246148" , x"8a6de4b1" , x"44e1667c" , x"deb47481" , x"db68b174" , x"43c88eeb" , x"5b095122" , x"516d4d70" , x"bf2c34bb" , x"1e84d803" , x"d8488020" , x"f098aa0e" , x"37966595" , x"a542e32c" , x"f7071b23" , x"7abe1a18" , x"b65241f9" , x"a3aa46bd" , x"fb901f13" , x"8b7283ce" , x"c288bdbe" , x"a5b63487" , x"3179830d" , x"8b3c1bc4" , x"5a434e63" , x"b89682f5" , x"3240bd3b" , x"85c24093" , x"d5026757" , x"fe636d0b" , x"f3dd402a" , x"37fb3118" , x"c4725d1c" , x"1b159878" , x"dca9fce6" , x"1c15220f" , x"74a660f2" , x"10478634" , x"552ac4a2" , x"67928dfe" , x"d6983478" , x"72c89121" , x"8de72e4b" , x"5da6210b" , x"1ef10bd2" , x"c3750a52" , x"3651ac43" , x"a0bdd13c" , x"7dc1db18" , x"c5a081b5" , x"68df2306" , x"eecf7dd5" , x"c26f5850" , x"f9058b66" , x"5b688fa4" , x"3128c503" , x"c593c55d" , x"238d4264" , x"fb463b64" , x"b23e82a1" , x"d89e0dfb" , x"180496cb" , x"d5a9c34a" , x"8680e729" , x"5e007521" , x"87c4a39b" , x"0cf5d266" , x"dc73a894" , x"f9be67af" , x"7c1f5901" , x"d7b3ee93" , x"64b98e4c" , x"de94f4bd" , x"abe2e950" , x"1353dd82" , x"bdc314aa" , x"0849cc4a" , x"8522289d" , x"9d2aa285" , x"5903b29b" , x"bc558b0f" , x"2666385d" , x"9d933aed" , x"960a212d" , x"a9a21ff8" , x"431bf48b" , x"f38610c1" , x"0b6157e8" , x"44113444" , x"c1434e70" , x"eb5cdceb" , x"3e272e6c" , x"1e4f3c74" , x"71414726" , x"502512f8" , x"b0136766" , x"df42f470" , x"5bf66147" , x"3bd012c2" , x"bc80c87d" , x"cedcebe7" , x"650b8c8d" , x"8e78dda9" , x"aef45791" , x"f18f4402" , x"b43c73df" , x"80f2b5cb" , x"713aed7a" , x"aa9a4b05" , x"05030a1c" , x"2728c323" , x"54b31a1a" , x"f925855f" , x"6c9f8c13" , x"a23e8c4c" , x"45307142" , x"2dbbfdff" , x"32721e2e" , x"12fb05d7" , x"d25c51c0" , x"7eb6aacd" , x"6e0f5443" , x"c935faad" , x"e344f51b" , x"76f54059" , x"64249192" , x"e20e5ce9" , x"c4e4ae3a" , x"a5b9f7db" , x"659420e6" , x"e73accd8" , x"cefac7bd" , x"01877c9f" , x"c14cbb80" , x"b18d4444" , x"609cfe97" , x"95c86f58" , x"374d0405" , x"1af8f529" , x"ca582092" , x"fd859ad0" , x"f30594c3" , x"3ae0c1e2" , x"53db540f" , x"553972a2" , x"abd7fb48" , x"b07b6500" , x"704b0980" , x"f61fab85" , x"d5604b93" , x"3a0265ee" , x"c4d3a1d4" , x"ec9b15b3" , x"2ad120d2" , x"e051ab9e" , x"dcaac0bf" , x"6e86cf38" , x"fd6842e6" , x"788c13c3" , x"83b14164" , x"8fe5f2b8" , x"e2603da2" , x"d66df6b1" , x"9688e031" , x"25f79219" , x"279dd996" , x"a3a7bc28" , x"332a35b5" , x"fedf3a56" , x"682e3122" , x"a3af54fb" , x"bfab2d85" , x"708445de" , x"d3597601" , x"0744757a" , x"ca3b0466" , x"154960a2" , x"518ace1f" , x"87c624d3" , x"88b86d2d" , x"c831404e" , x"170701f7" , x"bc94c80f" , x"1c98bf7b" , x"30ae63a0" , x"22e41189" , x"43071c8e" , x"adbc2855" , x"73c65029" , x"7ec3ebd0" , x"75c45269" , x"3090dc7e" , x"ac737bdb" , x"7eb8b3a1" , x"2d4ccbea" , x"25c9a708" , x"3015ae7f" , x"0e12c930" , x"18b35c18" , x"d9c84e4a" , x"52e9723d" , x"8f80d443" , x"2b9a8465" , x"edfad8cb" , x"0654f8e1" , x"b258c807" , x"d4a504c5" , x"9531c9f2" , x"3ead12af" , x"d0bddf2c" , x"245c67ff" , x"e1070e24" , x"27cb0b77" , x"fd294fc9" , x"4d921c60" , x"00223c00" , x"08983206" , x"dd8d6226" , x"68c7305d" , x"9cd127ee" , x"c87aca8d" , x"fd6d6067" , x"7180d254" , x"87160a9b" , x"047a1b7e" , x"7ac20b63" , x"49292a07" , x"cd251dc0" , x"f38ebbf4" , x"3a53ea35" , x"2bdb4d2a" , x"7f831b9e" , x"181a340d" , x"e69e44d6" , x"461f148f" , x"931cff63" , x"338c963f" , x"d85d98f4" , x"c0cc3bc3" , x"bd1787b8" , x"cd066f08" , x"96033f1d" , x"96099d00" , x"3f29fe61" , x"7f3b0868" , x"aa9a40d3" , x"974a05c7" , x"155f212f" , x"919c523d" , x"a03ee693" , x"2f62953a" , x"a933a98d" , x"e6d2f835" , x"bad10485" , x"064326b7" , x"e40854bd" , x"43ae2d36" , x"fb78395d" , x"c852eb99" , x"c4df1702" , x"998613fc" , x"94d9ad59" , x"8e642285" , x"eda5ecc0" , x"18b65ebc" , x"9480cd5b" , x"ed41ea5b" , x"0458fe6b" , x"65fcf92e" , x"1ef0a732" , x"0a371440" , x"dcda9c1d" , x"95ca3690" , x"7bfadb36" , x"69c8743b" , x"d848763a" , x"21291a12" , x"359b925b" , x"9be36cb7" , x"8d62f724" , x"0e2f1d68" , x"a1400984" , x"d929e929" , x"0830903e" , x"73ba7602" , x"9d5ddbce" , x"7c29e6fd" , x"5cc6ff75" , x"11443271" , x"0cae2adf" , x"3893d773" , x"7d547564" , x"a4f51632" , x"31485c61" , x"f9d01d4f" , x"1f826a8c" , x"f308198e" , x"349b440f" , x"bc89760f" , x"25820045" , x"6bbd0ff5" , x"306708b5" , x"af8c40a9" , x"0aeb44a5" , x"afabdb75" , x"a29c54bf" , x"3b344417" , x"48286d1a" , x"fea98ee7" , x"89e178c9" , x"6f83070f" , x"b1f6347d" , x"be6931ab" , x"7fc61130" , x"568a7ae6" , x"892a4212" , x"5ce80c3d" , x"71f78613" , x"fd68fd21" , x"1fba068e" , x"b99ebae3" , x"7d880e21" , x"d666d5ff" , x"da5e1640" , x"65e5a64b" , x"dfb9b4db" , x"da08bb6d" , x"4532027e" , x"2bee2b2c" , x"355db93f" , x"f2886e17" , x"90a28047" , x"59d45cd2" , x"a3eb79d5" , x"628767f7" , x"6ac268df" , x"6654b503" , x"34bacfae" , x"b7e6dcb7" , x"f2abbeba" , x"d5feb0f3" , x"15029e4d" , x"f36c7e94" , x"1b0fc5e8" , x"106116c3" , x"245cce9c" , x"aa1e5ac6" , x"2a9d26d7" , x"2d22c0b8" , x"9ef7254f" , x"5ef71ba3" , x"92dea4ac" , x"2b1c419c" , x"0d54fa1a" , x"1cfada02" , x"ee6336c4" , x"270f0d9a" , x"ba899262" , x"65409689" , x"bce330c8" , x"657f64dc" , x"103b470f" , x"0728ae6b" , x"dc45d525" , x"7335508f" , x"ef352c92" , x"193a2a5a" , x"fc01871e" , x"ea8024ad" , x"dbe36a04" , x"77608d53" , x"c91a64d5" , x"bfc6e79b" , x"836cb3d0" , x"bab552d8" , x"2d775ac2" , x"bc7e9caf" , x"6609f616" , x"a8138c73" , x"2249518c" , x"373ee1ff" , x"07e860a2" , x"0d2e9f40" , x"f06b9740" , x"0f06de19" , x"4d2264ed" , x"6be1514f" , x"4ba81ae2" , x"cf770e97" , x"553b4ff6" , x"511b0eee" , x"7791c7c8" , x"e253d494" , x"a5f054a6" , x"68bb4f55" , x"06755aa1" , x"3399e4ea" , x"d79ada44" , x"06872554" , x"8f1cc1d3" , x"11023da7" , x"daa64b53" , x"ad285725" , x"590e9c63" , x"14c15ce9" , x"722ecd7c" , x"54545077" , x"0de2a38c" , x"5e9cc7bc" , x"2d56eb5d" , x"cbfed9fe" , x"a9adca03" , x"2d2e229e" , x"54b13590" , x"17bbdf33" , x"e603301f" , x"0f42e5dc" , x"1e3f6b50" , x"4972b692" , x"fd08f50f" , x"b74ada18" , x"8a3c4458" , x"7e58c228" , x"b4f88a37" , x"e7b63daf" , x"ffdeaec9" , x"6790ca12" , x"49b07ea2" , x"113f92c9" , x"6a1e2620" , x"60019d8d" , x"76ffc013" , x"d93c71ed" , x"c392b0eb" , x"5d5d8276" , x"d175d1ff" , x"24822a91" , x"19a81e7e" , x"6bf48086" , x"2d991284" , x"de745487" , x"5c11089e" , x"ff3e1aec" , x"0e8432df" , x"88a01229" , x"859a4cb5" , x"65024cf6" , x"55fa32c3" , x"550f6841" , x"2cf8a548" , x"0b04217c" , x"357d8768" , x"db4496b7" , x"e7b824d1" , x"2e41e744" , x"ace66fb9" , x"55543535" , x"77ed882b" , x"6e6de4f5" , x"e981839f" , x"53d47730" , x"1aa080a4" , x"40a9c1d9" , x"bedc1b91" , x"21ae3f49" , x"bc7c0625" , x"172c6e63" , x"8fd6266d" , x"f3bfa71c" , x"2f275830" , x"4790391c" , x"98e2d7d3" , x"9402391d" , x"4cc8aba3" , x"5a5edcc0" , x"2255e170" , x"51247215" , x"366d0ddc" , x"c6d870ac" , x"e51ae5dd" , x"5ec415b2" , x"124abb52" , x"310541ec" , x"3e139975" , x"02d281c6" , x"0dc2d905" , x"646c19ac" , x"7114b24f" , x"e81bbe41" , x"03668716" , x"fcbe970f" , x"e5ae5507" , x"b57c01bc" , x"325830f8" , x"a350df89" , x"17e7214a" , x"9efd6dd4" , x"4eaf98cb" , x"ecd302cb" , x"74c031ec" , x"e178b217" , x"1a07016b" , x"04fad3ca" , x"fed1dc60" , x"b86c7970" , x"55040935" , x"9750cf8c" , x"4c1eebc5" , x"0e7783ce" , x"0fe2320f" , x"a386f8f1" , x"4c59b785" , x"4be58f35" , x"0bddad32" , x"76ed671d" , x"8163bd16" , x"f2abc08a" , x"c2ecce9d" , x"8d4b720c" , x"a18dcda5" , x"80df7f8f" , x"170323bb" , x"222256de" , x"14b3664f" , x"b68f620f" , x"c6f93c4c" , x"ecd35ca7" , x"e7b6e901" , x"e74ef9ad" , x"88a54754" , x"a2e40e63" , x"1bf187ca" , x"578b485f" , x"d3683585" , x"a9e52fec" , x"568d927d" , x"a8dc3a09" , x"4b41d16e" , x"453b707e" , x"bf0e658a" , x"a46c783f" , x"02a56ba2" , x"6de39386" , x"0c670b73" , x"cd5dcf9b" , x"aafc8d1a" , x"5509fb61" , x"9a7ce0ab" , x"b5e3c317" , x"86aea6b7" , x"a77ec27a" , x"bace3d0c" , x"3d9b957c" , x"b50e9075" , x"eb4b4481" , x"c8085396" , x"9a9514e0" , x"49b8dbf9" , x"621c603a" , x"b149c6b1" , x"c7b64df4" , x"8e81ea1d" , x"7eb8a175" , x"658262f3" , x"e2935501" , x"0fc467e4" , x"65e283f7" , x"c7b99565" , x"4726ee02" , x"566be57d" , x"3e16356e" , x"9b9d19b7" , x"0061bbbe" , x"bdc2d35a" , x"651de231" , x"1ad50a77" , x"33b61972" , x"20bd4af2" , x"c5a6b0fe" , x"8caea916" , x"9bc3d23a" , x"7c37fe8e" , x"c7704699" , x"e3f636db" , x"7fd82ae7" , x"cc88a93d" , x"626f5384" , x"bbfdc6e4" , x"d4aac7fd" , x"0d241625" , x"20c1cd84" , x"12a89c78" , x"3fea0c3e" , x"16a9bc57" , x"80ce9bdd" , x"cc60b8e6" , x"20d276cb" , x"f168fb2c" , x"fa8b34eb" , x"af07fbcd" , x"ba141b80" , x"21d0304c" , x"3930ada6" , x"b90479a1" , x"aebd5e13" , x"1c40202e" , x"72de8777" , x"1e1402f2" , x"ac0c0dc2" , x"a40616f0" , x"e8cc2e4f" , x"542d2b18" , x"d6b91d93" , x"a760399f" , x"363e6252" , x"bfc71451" , x"f37955b9" , x"954ba8e0" , x"e0bd814c" , x"bd72c22d" , x"b585a23a" , x"3c1d9dc8" , x"f880ac8a" , x"bc262d6c" , x"6c43ca6e" , x"f8792500" , x"d657bf17" , x"ddef24cb" , x"17e3c607" , x"16137752" , x"ac65b025" , x"5dceca5b" , x"192ed0ed" , x"5e83d012" , x"b28ecf43" , x"af5e06bd" , x"374895e4" , x"9912b3fd" , x"c71fde34" , x"ca13c16e" , x"14ab277d" , x"5e1e8061" , x"67c1d12f" , x"34be3de4" , x"351e17ed" , x"162fc765" , x"15c4b379" , x"c59d7614" , x"84e92585" , x"34a715cb" , x"fa7e24ee" , x"6365c519" , x"2a84e35f" , x"8d415b88" , x"eb2124bc" , x"3a9cae21" , x"4e043871" , x"a456387e" , x"94b52a84" , x"7c06e7c7" , x"d8085e5f" , x"26df592b" , x"6358b3f9" , x"c82cb19c" , x"018a1a7f" , x"19c15612" , x"028a1af1" , x"4b47ee7c" , x"32c88faf" , x"3cc47a70" , x"64b4b01a" , x"87e73e85" , x"324f2c6e" , x"176c75fc" , x"d5d37d33" , x"67c2c057" , x"c79cf98b" , x"1ad73437" , x"13c39a23" , x"1cbea45c" , x"4a9a7e53" , x"c8d04433" , x"4685deff" , x"4aa45a27" , x"9f281fb6" , x"9a812ade" , x"ebd1e00f" , x"f6e4676c" , x"39b5049d" , x"6eb75633" , x"48e85c91" , x"b1db47b4" , x"15aa8ed3" , x"c212cb53" , x"53ea8253" , x"6ec1a5cf" , x"0d565978" , x"a7ceb820" , x"9c62ead7" , x"1c18e837" , x"8b691ea8" , x"ef0ae2b2" , x"5910390c" , x"2ffd6e67" , x"86e7481c" , x"44244bde" , x"fff6e8f1" , x"cc3e9a8d" , x"daf19f53" , x"7cd399c0" , x"e7289cea" , x"c4da72e4" , x"20f9655b" , x"6560b2b8" , x"9da640d1" , x"45df5103" , x"d49142d0" , x"0988357a" , x"fce27b2c" , x"ac5d0e24" , x"a5474262" , x"6df7efbb" , x"c015c711" , x"73a52eaa" , x"c1e3203f" , x"9c1f996a" , x"aaa93160" , x"0f350df4" , x"8a3f3e0d" , x"50d904b0" , x"baf1f8f2" , x"c5d11e0e" , x"c79d2874" , x"b2496eb7" , x"7d17f8d5" , x"2015c514" , x"9800916d" , x"21519ae5" , x"f798a8f2" , x"17a4672d" , x"14108f18" , x"020082d2" , x"0900d865" , x"6c50e584" , x"5f493e14" , x"a7d3a4da" , x"13f22216" , x"b9117347" , x"c8c0818f" , x"87fd551c" , x"7a2487e2" , x"1bdb7e09" , x"70ce9889" , x"a1bb70f6" , x"48239825" , x"20624b99" , x"844d5547" , x"2261b391" , x"5e2c1cac" , x"193d7667" , x"1e2e22f6" , x"245be5c1" , x"993f7cda" , x"2b128462" , x"043ec379" , x"323d5e92" , x"77c03ecc" , x"51465aca" , x"1b441d0d" , x"51017db1" , x"56b6f38e" , x"37b23aa1" , x"163e8d8f" , x"4044474c" , x"34853b65" , x"e4969009" , x"848d2a8c" , x"b4066fe1" , x"7a0e33b6" , x"8e44d787" , x"090239e1" , x"2f370b6e" , x"da675280" , x"3647a734" , x"f35b6e15" , x"13cd0012" , x"da59fa7c" , x"e9eed2d0" , x"faf4f631" , x"b4eb49c1" , x"dcc02ddc" , x"8ecb41ee" , x"d2412d51" , x"503ce1c1" , x"eb2af3ff" , x"2a8c511e" , x"9925b74c" , x"9f5bfae1" , x"d3a77d84" , x"fce94a64" , x"89a08e3c" , x"2ba16ec6" , x"e9c371f3" , x"41feac41" , x"2af3c7fa" , x"6594a3e7" , x"04d5e266" , x"12f1523a" , x"db4397cb" , x"af20eb6a" , x"d76476e2" , x"6702ebf4" , x"c9c69f17" , x"fb9b1675" , x"bac1ba06" , x"66f58780" , x"bc0b4da9" , x"9ee45b58" , x"962276e7" , x"2784c798" , x"902fd5ac" , x"619fd6da" , x"ec9a80c4" , x"29401365" , x"9af0d2db" , x"c213a805" , x"19f03fa3" , x"df01237f" , x"9e77bce4" , x"59cc8126" , x"bbdba2c9" , x"af7f44a8" , x"4a7ca0e0" , x"4b4d532e" , x"51916628" , x"87d7527f" , x"92eaa3ca" , x"d519b2f1" , x"a429dc54" , x"98f51e10" , x"0e301d60" , x"55d6f69e" , x"fadbb1fb" , x"4c9a02c8" , x"cae25d94" , x"73dd1ac7" , x"a3a150ff" , x"6c328167" , x"53070d6e" , x"5c0f28cf" , x"f9017e68" , x"8eee01c7" , x"81571412" , x"be1773e9" , x"ebe3b6f7" , x"6ca1345b" , x"91d2145a" , x"6dea42c2" , x"7243c56a" , x"1ff7a935" , x"f6e735ba" , x"06414ec1" , x"1ec536ac" , x"4a4994c0" , x"fc23f7f6" , x"51490760" , x"3adf4d48" , x"a7583c9b" , x"98d4b9a9" , x"f4f9c0ab" , x"92024f3e" , x"ef8c0ee4" , x"c3bfb04f" , x"753809fe" , x"6984ccb2" , x"3d8ffe15" , x"0e4e7760" , x"c38ed0c1" , x"818953f4" , x"c2634781" , x"2c0ae592" , x"bd9b1c94" , x"876e3f07" , x"be625be6" , x"88d61be0" , x"1b1d99a9" , x"aec470e3" , x"ae7abe82" , x"78f1065d" , x"76983ecc" , x"54b0410c" , x"365053e1" , x"5fe0365d" , x"1938863b" , x"234f1c62" , x"d2d5c6d9" , x"bab9490b" , x"2ccd7029" , x"544cf732" , x"29dfb7a6" , x"a916f8bc" , x"aa7e2376" , x"10517fc4" , x"e4f6b3a9" , x"e84a6d7a" , x"843d28ad" , x"1acae058" , x"b3e44c7a" , x"19688a51" , x"2751b2f8" , x"647c34b3" , x"f415c320" , x"aa694f1e" , x"8a77610d" , x"7edf8973" , x"ae030a7e" , x"765f54d0" , x"095c31a1" , x"3616dcb8" , x"cf27fbd6" , x"68d52d36" , x"bfa57c96" , x"1b93d549" , x"1ec49391" , x"7d4425d4" , x"86695c39" , x"1ca06ed6" , x"5369d527" , x"5bcd20c6" , x"8be41c5c" , x"4a68d9c3" , x"661d0c8d" , x"53eaef35" , x"6a438f62" , x"424fb511" , x"2e44d46f" , x"8b92b330" , x"41610693" , x"11d3638a" , x"0541d53f" , x"04707e4b" , x"ec760158" , x"228a1066" , x"a758e029" , x"e583a350" , x"eebfc341" , x"be08da53" , x"29dbf25c" , x"9a89abf7" , x"ebcd0799" , x"f3f04ba6" , x"cb6eb2fe" , x"ea069391" , x"93d01b24" , x"3e0abf05" , x"70a62c38" , x"e6ede86a" , x"41f2f950" , x"717133d1" , x"c07f8f0e" , x"900bf22e" , x"3a8a155c" , x"59e41e60" , x"106e90b0" , x"0963bc2f" , x"c46fb4e8" , x"90541acd" , x"abd3e80c" , x"58e16226" , x"b7182aca" , x"c58f9082" , x"a45e1929" , x"a1541882" , x"6b46bfb4" , x"e48200ee" , x"6408fbd0" , x"dcab9be7" , x"d0ee8ece" , x"566dbeca" , x"5142f3cf" , x"a9ed9c83" , x"d085ada0" , x"af324efc" , x"ca00b8d5" , x"666bb61a" , x"da2df775" , x"04b55856" , x"817166c9" , x"010bc7b3" , x"a2bab478" , x"63ea9a9a" , x"f36dd0eb" , x"fffc2bd5" , x"71a7a299" , x"33376ddf" , x"0f5d64be" , x"a0c76885" , x"dde35221" , x"eb6335d3" , x"a19595bd" , x"da4ff304" , x"5ae61b4f" , x"d3ed74d8" , x"ff3b9b30" , x"ec71c819" , x"39634da8" , x"469f649c" , x"a707088c" , x"a51f5b76" , x"9ae0aaba" , x"6b0e612b" , x"6322842e" , x"fdf6bac0" , x"246660a7" , x"7882c7d4" , x"066f3f17" , x"ace2d0e7" , x"6bce032b" , x"eeeeb979" , x"2f213246" , x"9233ce13" , x"b9cc687c" , x"703733ba" , x"5ed016cb" , x"51ee8b31" , x"d7707b46" , x"ea5bd791" , x"bbf67a05" , x"fb6b6fcf" , x"922ec070" , x"479ac0a2" , x"2d465f93" , x"05101e8b" , x"f5171e9f" , x"5617ab37" , x"43ec2503" , x"e2da9003" , x"ecb15570" , x"1c7be16c" , x"3949047b" , x"4fe44d8c" , x"5fa1e0b9" , x"865aebcd" , x"16666c57" , x"1e8f5de9" , x"a3dead8e" , x"c2c8cd0f" , x"2e3ce889" , x"500a0ae9" , x"0b887832" , x"49fb0cac" , x"b921e5a5" , x"53684e81" , x"58f1ac65" , x"69625c78" , x"a91e2f26" , x"436b3301" , x"6245367e" , x"7c85ea07" , x"a099c7c1" , x"3a09933c" , x"058ad79a" , x"ee69bc61" , x"e91b1d72" , x"0b676e23" , x"ccf1697a" , x"f9fa436c" , x"beefdc5e" , x"c8726697" , x"d0282955" , x"735586ec" , x"62205cec" , x"36c6413a" , x"9e060308" , x"1a64a160" , x"9353a181" , x"8b847e72" , x"87b177e7" , x"893d0273" , x"466af8a4" , x"aafdc83b" , x"3fa625d1" , x"14b17e29" , x"739e9922" , x"a59332da" , x"3a4b6351" , x"254f6141" , x"cdf0686e" , x"67310e80" , x"fc7153d5" , x"eb1eda59" , x"07ad8d65" , x"6c66fd97" , x"892149cb" , x"a46ec92a" , x"164ab140" , x"9d9b82fb" , x"cd55dd49" , x"ccb5ab98" , x"fd3899c0" , x"7157b906" , x"112363df" , x"b3436262" , x"f07c692d" , x"d1ae2ee0" , x"04a74860" , x"43eeb0da" , x"af100c24" , x"0e42b551" , x"c8a2f426" , x"b51ddbf5" , x"88bd3d50" , x"ccf86b3e" , x"e2a6eaa2" , x"f7a1528b" , x"e6252f59" , x"fdf71ba0" , x"a03d72c1" , x"0ad01711" , x"234b61cb" , x"ec5af39a" , x"37c1d87e" , x"1015004e" , x"2ea0cc20" , x"61a94d4c" , x"0ab4b4f6" , x"20b23117" , x"1b608754" , x"706cd381" , x"9dcf3d8f" , x"0233c6f9" , x"f08d9fa2" , x"dfbeae3f" , x"5abd9c4d" , x"e3135b87" , x"691efce3" , x"84bc1ca1" , x"fbfe52c9" , x"4e477293" , x"f2117a59" , x"657a2c5d" , x"ad3895ec" , x"67136e10" , x"fd016092" , x"39964727" , x"c44f0fcc" , x"8d21f76f" , x"5631ec59" , x"49306e03" , x"a991db89" , x"5f0907dd" , x"3e819dd3" , x"0ca9643e" , x"4ba65cfa" , x"d06badb5" , x"ae202b6a" , x"9f0d6c09" , x"8720f852" , x"4f9165c8" , x"695e314e" , x"3aa61704" , x"9a467f8b" , x"6e49d108" , x"c0221507" , x"b979edd0" , x"95626e10" , x"dcb07ff6" , x"8d424628" , x"ae9ede39" , x"9564e24c" , x"93c4565d" , x"8306a14f" , x"cd4dcd33" , x"1524cc0a" , x"2ac663cd" , x"b835bf9c" , x"a332d3f4" , x"ff04163b" , x"fdd83fd0" , x"5ac2c28b" , x"e8ccf1a1" , x"f8a46af9" , x"7950c3f4" , x"58b0ddb1" , x"9c32b2f7" , x"e2f489d4" , x"e5d72a24" , x"7466e1ee" , x"b665212d" , x"69d65eeb" , x"6cf25d12" , x"37bd49f4" , x"871490cc" , x"202ae62e" , x"3a84d2b8" , x"4f1506c1" , x"e50348d9" , x"b9e1faeb" , x"1bd95560" , x"c86a4dc2" , x"f32d2d80" , x"b19c10a2" , x"65e893f6" , x"02826688" , x"072d0b3f" , x"d7dcd444" , x"7272f590" , x"ec1df337" , x"34b6fc63" , x"c55d4161" , x"e40fb6d2" , x"0aebc191" , x"f0beae67" , x"60d0ce95" , x"13733aa0" , x"b44f9a00" , x"2376c0fc" , x"bac15dee" , x"839521e3" , x"396a38cf" , x"ddf962fc" , x"44e0c54e" , x"ce67bdf6" , x"ac4bc52d" , x"d70d4086" , x"7a3cedb8" , x"eaa801cb" , x"9fabe0ea" , x"d314b265" , x"3c87a7ab" , x"a7fb2732" , x"2d57fb70" , x"e751ecd5" , x"d4638254" , x"474f8b57" , x"c454fa7a" , x"d3018121" , x"ef39f7c1" , x"aeec97c4" , x"1b9e9b60" , x"b7823b4e" , x"2ea6762c" , x"c7e7d0c4" , x"195e4ee5" , x"a989eb1d" , x"7d612906" , x"c034e4b8" , x"317886b7" , x"33bf82ef" , x"e5592669" , x"919bc0c1" , x"195df06b" , x"a60b3eba" , x"0b4e6f4a" , x"b2a35ec4" , x"8eaae525" , x"a3349626" , x"c5c23c8d" , x"cf23293f" , x"4fdb4da2" , x"ca1217c2" , x"2dd1cbb6" , x"b9b24fa8" , x"56c5cca6" , x"06f088da" , x"35cc1aae" , x"f3fe3e73" , x"82995b06" , x"22e8f255" , x"e8077e17" , x"357b6ea0" , x"a10128dc" , x"217739d5" , x"19fe1ff3" , x"df139f6b" , x"640f0e97" , x"e3911f11" , x"0dfb5adf" , x"01a16f0f" , x"805413b6" , x"b202e6ac" , x"6e85475c" , x"d1de7cf5" , x"ff601d6d" , x"a7878a40" , x"cfc52fc9" , x"75caf69e" , x"7c53aae4" , x"bbad9deb" , x"e4fa872c" , x"9123f46a" , x"233640f9" , x"719b0cc0" , x"63d75cbc" , x"869300ff" , x"ed6737a5" , x"90df28bb" , x"eae0e02b" , x"a4124873" , x"b6acc95f" , x"9895bb6d" , x"9e4b5bc2" , x"c4674c7c" , x"57e1b718" , x"ad9867ae" , x"ef9f7cbd" , x"225be46f" , x"1ff1310f" , x"403674c3" , x"bb07a479" , x"54d3a8db" , x"a57f8b99" , x"2ef7a531" , x"d54972d5" , x"98606d22" , x"65f5d2e4" , x"c638a025" , x"bff4593e" , x"5825ad31" , x"d5d102e5" , x"4b9db004" , x"528cc3b5" , x"e76896d0" , x"8d61047c" , x"79f11591" , x"faa834f2" , x"92ea54f8" , x"8c9f7be6" , x"45d19b01" , x"5496a458" , x"28b16b5f" , x"9e95b019" , x"b2539ba7" , x"5c52ada5" , x"31917eed" , x"c1aa9c10" , x"239f3650" , x"69f5665a" , x"1b5071d8" , x"7e0a5431" , x"4d6e9edc" , x"b1dab156" , x"4b5ffa5e" , x"f905168c" , x"0107916c" , x"53e7bfd6" , x"235e1d66" , x"d67a44f1" , x"be751c65" , x"bd33d662" , x"2c2c67df" , x"f444c6f6" , x"a6a13630" , x"082c14de" , x"cdc679c0" , x"5b5bc40c" , x"84e2b396" , x"a9a3ae9c" , x"16a924e3" , x"48107c6b" , x"b286b612" , x"3afa6277" , x"dd7204d3" , x"b60c854a" , x"749224bb" , x"9fe402a9" , x"e3a0f034" , x"973220e5" , x"883213b9" , x"a9127665" , x"52cb8521" , x"0c2c8b1f" , x"2e5e42b0" , x"5949f600" , x"8f237ba2" , x"738b0e70" , x"3fe27659" , x"3dabf323" , x"60973e9f" , x"b70d30b4" , x"1a332012" , x"db2ec337" , x"fca68fdf" , x"4810e379" , x"40da2a07" , x"bb2625a6" , x"6b045f0b" , x"23446dc7" , x"6fca1bef" , x"d63376c1" , x"bb77285f" , x"237b66f7" , x"62436e29" , x"9694e3e7" , x"4b95c832" , x"5dbc73b8" , x"d94bafa9" , x"ce87cb2f" , x"2071414d" , x"80f7c703" , x"7a181bfc" , x"7d560df3" , x"c8fd096c" , x"e08643c0" , x"ff7f9eb4" , x"5a678073" , x"cb623af1" , x"730ebbb9" , x"06fd1a16" , x"f6a9ebb6" , x"f5958a6d" , x"0ad40741" , x"55e2dfe5" , x"f913cc2a" , x"0c098e92" , x"306fdc0f" , x"9b1ebc77" , x"aac86546" , x"f95bcf9a" , x"9620e80a" , x"b0ff9409" , x"acd42ada" , x"acab0448" , x"5c6bf0e0" , x"336863de" , x"9eca9125" , x"357a2119" , x"cfa79581" , x"dd047645" , x"04ee0ede" , x"dd93db8f" , x"1578bbe7" , x"b89b520d" , x"f98c9a32" , x"0529bd60" , x"a6bed7d2" , x"5fe9220c" , x"3b3266c6" , x"5031e030" , x"674b320f" , x"7f90ef75" , x"1f3cbc8d" , x"baabc2c5" , x"44b8681c" , x"b70661c8" , x"420234f7" , x"20428a16" , x"54e8034b" , x"ccf4fe02" , x"26f8cefe" , x"54ae7c8b" , x"591707b5" , x"69e7d7a4" , x"1f25023e" , x"5444cd23" , x"e257daca" , x"9d8ba71f" , x"1822a0e2" , x"505c3d77" , x"ee172475" , x"c8aa0b7d" , x"66262c22" , x"aba28198" , x"0c22809f" , x"89951216" , x"57a5ca39" , x"b8bd1796" , x"bc684722" , x"bad30960" , x"cb704a2a" , x"a3b515aa" , x"8b7ef3fe" , x"a2ddf00f" , x"afac574a" , x"1a1d5519" , x"e4c51cd2" , x"1d5e7a17" , x"0e06d5a8" , x"8e5b3ed3" , x"4dbcc089" , x"778ae5ee" , x"0bd335ac" , x"be5cdb35" , x"320ac3e1" , x"177b0e82" , x"b85cc92e" , x"cc0c6fb7" , x"b8c4d288" , x"8baef279" , x"e0b7709f" , x"f8709ced" , x"951a53a7" , x"34afa17c" , x"12185e55" , x"e699ec0c" , x"ec38fcf8" , x"bc30980b" , x"cce52f6e" , x"ca3b9729" , x"4933d034" , x"65c1786d" , x"8b2d8366" , x"e8baf276" , x"fc1a4bbb" , x"1d556ec4" , x"b736ad8d" , x"262fc8de" , x"d6c6b637" , x"36f7123e" , x"6eea2a11" , x"2167f02b" , x"787adc86" , x"11c1517d" , x"8f8aea1e" , x"16eb7779" , x"44e32ee3" , x"98c43010" , x"bfbfac9c" , x"f4fa4075" , x"80feca0b" , x"1eefbaff" , x"a595516e" , x"db06b095" , x"4ec86a02" , x"d27db2b8" , x"23837536" , x"78d74fc2" , x"79bf25da" , x"ac2fbb0a" , x"5cca21a2" , x"29fc4d57" , x"c9c1cd34" , x"c414e2c9" , x"c7c17796" , x"3dd8efd7" , x"ab239dc4" , x"89906d14" , x"222d4f06" , x"b914b4b5" , x"0584afc7" , x"349a2eda" , x"8f51b879" , x"95892f34" , x"4d0279aa" , x"24fc7eca" , x"f07d27b1" , x"750cbd8b" , x"fb1c8026" , x"6aca3bb5" , x"495ff422" , x"65575686" , x"cd028ef7" , x"73710096" , x"e5678dbe" , x"9fd1b530" , x"98f7806f" , x"8f6324dc" , x"e24eeba1" , x"c8676293" , x"f19863f6" , x"4d1de71a" , x"8c959fd3" , x"ce6b4c17" , x"ba778f08" , x"b3c2a9fc" , x"93a66e87" , x"57f96772" , x"069e9871" , x"05465986" , x"724fdab2" , x"6312c49c" , x"a5740b9a" , x"514b7948" , x"856d8e8e" , x"227410a0" , x"5f4fe1ea" , x"6f7a5c51" , x"efe80ead" , x"bf143d23" , x"d45c436e" , x"02662bda" , x"d95daa60" , x"ff4d8388" , x"5f5e676f" , x"4811e68f" , x"97daf1ba" , x"f870c7af" , x"df5f9ad6" , x"c99e15de" , x"eef9f614" , x"fa694b2f" , x"ab207991" , x"27696e0c" , x"34ef4d57" , x"634fdd2c" , x"a762c08f" , x"eb084d11" , x"1271f868" , x"80f33888" , x"681f414f" , x"75b1bd04" , x"aabc0664" , x"1e60f64c" , x"ef08a51f" , x"997c83df" , x"cf9a6bc4" , x"d93a5b53" , x"7c0b5b15" , x"26eab470" , x"c1ba50e5" , x"a40aab3c" , x"6ac39f39" , x"b5a45ded" , x"f8c6f782" , x"14cc9a3d" , x"fcebe8fb" , x"b87e8e2a" , x"dd38c5c5" , x"00dda5ea" , x"638de300" , x"dbe93654" , x"7469f5c1" , x"fc68f121" , x"3f26e470" , x"31945ad9" , x"c8cff3b3" , x"5620c800" , x"e201a538" , x"9d43e80e" , x"e9e9023d" , x"e903750e" , x"8eebc2c0" , x"0675d1f6" , x"994f6b8e" , x"1f4cd75a" , x"261cc8f9" , x"27e253f2" , x"e6539f66" , x"becf4148" , x"734cfe61" , x"19d559be" , x"34a6f158" , x"1d842a32" , x"e64f86e5" , x"f067712a" , x"c338ce50" , x"801590f8" , x"e1ea9f69" , x"2b9ddd8c" , x"48f27f54" , x"db3cc749" , x"ac5889d8" , x"5509cd68" , x"aa0e3f66" , x"86ec9d32" , x"1f70cdb6" , x"720e2342" , x"68460523" , x"50b2cc69" , x"467934af" , x"2754dae3" , x"b777ab07" , x"509f9247" , x"488be0e7" , x"da59043d" , x"e56d49c3" , x"670ca230" , x"d39aac9b" , x"f067b9a7" , x"63d8c707" , x"68df5306" , x"7f769128" , x"c4e81c25" , x"b1dec0d1" , x"5cf468b3" , x"d59934fd" , x"a429d26f" , x"9c10b0fd" , x"de9f89ee" , x"9321f971" , x"ed64b019" , x"53777ffc" , x"69d78350" , x"74d83e14" , x"edfc1fa0" , x"b6bb4eba" , x"701fdd6d" , x"e2685e79" , x"cf05bac9" , x"b889ff5b" , x"5a5be0fa" , x"04c3ce8f" , x"55e6b1c6" , x"acbe2683" , x"536947d0" , x"70421d41" , x"18d36cc6" , x"7014fbb7" , x"b86248d3" , x"1df62005" , x"01a32245" , x"d08efaa3" , x"690f06bf" , x"5329b9c8" , x"e6c423cd" , x"3f08ce45" , x"0ff2c3b8" , x"57bc0dbc" , x"e50ce83a" , x"602d5c20" , x"75a4bb03" , x"8beaf300" , x"565e548a" , x"8fd9ffc4" , x"6c49006c" , x"65549b00" , x"37c2650a" , x"65ebe7d3" , x"18eb1e32" , x"83ef1b22" , x"3f8da73e" , x"a853ebed" , x"73627ca0" , x"f36f2db5" , x"6e89f1fe" , x"b8ebd50d" , x"6ace6b9b" , x"666ba04b" , x"70fc6976" , x"d4f58535" , x"2735c3c9" , x"2263ff60" , x"0296e262" , x"0f7ac01b" , x"bfcf5e0a" , x"159136e7" , x"f3ce91d4" , x"29f53d7e" , x"e8c39289" , x"530013aa" , x"12ff51a4" , x"4d3df757" , x"835f1a89" , x"02fd8691" , x"171e0df3" , x"8a37386a" , x"08393eb7" , x"186a584d" , x"1e24c526" , x"2581ff69" , x"266151ee" , x"a1927847" , x"da4c2e72" , x"dbfc6c3b" , x"3ef9a58b" , x"f96696b0" , x"e9cef112" , x"92227788" , x"ca5842c9" , x"ff319347" , x"f4e140c5" , x"8db4e684" , x"591e1765" , x"83f515cc" , x"afe31ba4" , x"54a7947a" , x"966a5055" , x"6e149911" , x"6a910ba6" , x"7de703b5" , x"f992286d" , x"122f7c99" , x"01acba73" , x"e342e09e" , x"90b7ba7c" , x"108bd3af" , x"be4aca2e" , x"6fa9d12e" , x"befd7fb0" , x"d39dfdc8" , x"46b1ad06" , x"65003992" , x"ef593901" , x"9d0cb098" , x"cebb8891" , x"d192706a" , x"82cfd92d" , x"e2e04ca2" , x"6abed3fd" , x"ee5d54f7" , x"27dd1397" , x"30d7433f" , x"fe39732a" , x"42327256" , x"495b7f8e" , x"e5da8691" , x"44b7c36d" , x"97e6901f" , x"c86a9c55" , x"80fba9f1" , x"0f91c44c" , x"9ce116d6" , x"b5ca9d96" , x"d1c5a7fe" , x"a001d676" , x"8829e375" , x"e08cbb9d" , x"33bb3190" , x"5817aac6" , x"74325cbf" , x"b7ba3eed" , x"6d8b91fa" , x"71d4cff6" , x"f74f3bbe" , x"2e5af513" , x"9ebbed9a" , x"99c84083" , x"b2051378" , x"6ba38233" , x"b85cb54d" , x"02d47b19" , x"58ce1f87" , x"4b66652b" , x"84597be9" , x"a4030f9f" , x"8e838a1b" , x"b2ce4cef" , x"28101216" , x"c099f5bd" , x"8fe2e7aa" , x"71a7bfe5" , x"b1dea0d0" , x"defe0f4f" , x"6d2c30b7" , x"1896cb67" , x"d615d16b" , x"db55e007" , x"bb3c2ecf" , x"4f102904" , x"5c2afe97" , x"7a6cee4e" , x"7447431c" , x"9464399b" , x"62ea72ce" , x"4faa4393" , x"c68abfc1" , x"05d0f501" , x"bbf930fb" , x"8a8d0b6a" , x"6e26b042" , x"c64b79ab" , x"b199c4c3" , x"4b5e2792" , x"f1f982d9" , x"b90362aa" , x"c8c377ae" , x"8ee64411" , x"b4a05b6d" , x"bd350709" , x"1bfd5424" , x"38b88434" , x"63d27ecb" , x"e18f2357" , x"97458845" , x"61241470" , x"7599ee43" , x"539a2bc4" , x"0ce314c5" , x"a5cc8ee4" , x"3a8b44eb" , x"f2f1defe" , x"d58d6a19" , x"7f5cd65f" , x"04014a6e" , x"1be682bd" , x"dd1c27b0" , x"f4eb22de" , x"13fc554f" , x"ecd4fb7c" , x"ab466007" , x"6040564b" , x"800dd978" , x"77026d80" , x"37ce7111" , x"62e6d76a" , x"9255687b" , x"f3eb45c9" , x"1f47c9d4" , x"39230375" , x"abd18cd2" , x"e6ed1eae" , x"997e7043" , x"02bbd7bd" , x"0e547419" , x"aab0c2d6" , x"0e6c7ee1" , x"f0035b7e" , x"270a482d" , x"045bb460" , x"0505e2e4" , x"00910812" , x"6f67aa24" , x"064c8450" , x"d50c7779" , x"9af2d732" , x"9e0d4842" , x"1a231262" , x"85273399" , x"6393f1d9" , x"dd2677d3" , x"2c6d8ec1" , x"1902bb1f" , x"9b201e55" , x"e8761be6" , x"9dfbbdce" , x"1ba6fb7b" , x"45ea5267" , x"8459e65e" , x"4150b1dc" , x"24a5df99" , x"08986603" , x"8f32e8f4" , x"56868ec3" , x"012c2154" , x"b8a763b3" , x"c4454561" , x"f416f30d" , x"d9450218" , x"1b9d3f4a" , x"eab4cc6d" , x"e022c7fa" , x"fca9f3f8" , x"7315341e" , x"81506727" , x"42d2e804" , x"457be328" , x"c26743f8" , x"19cac905" , x"ce0e43f5" , x"82026188" , x"3dcc2da9" , x"95ea7ad1" , x"59079ed5" , x"c34c9198" , x"bbd0fe56" , x"153d0a42" , x"45c12572" , x"a95e5e3c" , x"e3963d79" , x"8458bc86" , x"c70d49c4" , x"2bc9cd9d" , x"4a8a1922" , x"f0455409" , x"25abc32c" , x"9729e7da" , x"7552fc44" , x"70cd6f33" , x"bacf46bf" , x"f121995d" , x"c95cb308" , x"a7e9f7cc" , x"b7fda22c" , x"73b2b6c8" , x"46ba203d" , x"d6f66900" , x"04365608" , x"885a0392" , x"61aa956c" , x"8dcb8afd" , x"8a01e5d9" , x"ae18c64e" , x"56c26f09" , x"5e002853" , x"d6134fe0" , x"3d422633" , x"7ebaf78d" , x"94345463" , x"d7fbb830" , x"ddec4f4d" , x"e9274abe" , x"68228590" , x"8f2d85d5" , x"1cd45884" , x"5de5625d" , x"719fe176" , x"c9aa0f8c" , x"4cd8e28d" , x"4fdd45ff" , x"66c149fc" , x"916baef6" , x"d5575093" , x"15ac8268" , x"6754355a" , x"12ba1279" , x"63e291e0" , x"efa816c6" , x"5c4660e4" , x"87892170" , x"23e7c671" , x"a9353c67" , x"4297e460" , x"a3520c22" , x"163983b4" , x"98243e7a" , x"6decfbc6" , x"fe2f2613" , x"41dd48cc" , x"d3486877" , x"4c2c96f0" , x"9d6c12c2" , x"6cc38541" , x"bd9d6ec6" , x"1e845dfe" , x"85481f55" , x"7ebcb4a8" , x"b86f32da" , x"b4d71ab7" , x"1f746f7c" , x"3e5ad30f" , x"aeba94b3" , x"c8fa5a47" , x"b7cbf943" , x"12f788c0" , x"acbcbe1a" , x"64d58b5a" , x"aa951393" , x"00de6fea" , x"790adc59" , x"387e47e6" , x"0eae9f19" , x"00553bf7" , x"60483763" , x"306e1421" , x"9fec657f" , x"2479d5d3" , x"1d42a654" , x"44a0a0e3" , x"889e90fc" , x"2cc5b9ea" , x"a793a03a" , x"237e7fbc" , x"f4e9f14f" , x"9950913e" , x"f4998ea1" , x"e6abbb09" , x"e5ad2d4c" , x"f07b3130" , x"e7f9bb88" , x"389f8b7f" , x"25229883" , x"7b9059f9" , x"6057ef1c" , x"604243b0" , x"aea260a6" , x"861672cb" , x"88875552" , x"43ceb0a3" , x"b72ee312" , x"117fdbd4" , x"d2f0fe8c" , x"6fb321b0" , x"01172405" , x"2c81a1fa" , x"ae57f3fd" , x"06aef49c" , x"bdbf63a2" , x"f465cb88" , x"eb049e7e" , x"6e3b92c6" , x"948a782e" , x"f628b3e5" , x"055969dc" , x"c32d986e" , x"d6510a20" , x"01e19a1f" , x"98d952c6" , x"ae170325" , x"46573ddf" , x"b4b9305c" , x"50af1430" , x"a5272913" , x"017eb639" , x"8d642d9a" , x"7b5b3a86" , x"37d5f940" , x"2b215c18" , x"c5b9cac4" , x"6006e5d6" , x"3a601079" , x"8367b551" , x"5ef0fd6f" , x"f9d919e1" , x"e413e945" , x"2af41d90" , x"db3b844c" , x"ddf09e6c" , x"6705e285" , x"ba186e84" , x"5169b372" , x"6935c73e" , x"9bcf881c" , x"ae1cfe4a" , x"e9028deb" , x"5d065c14" , x"e8baa8b6" , x"4ba9474d" , x"9772bb29" , x"7607fb26" , x"55236652" , x"b0ba22d0" , x"da6260cb" , x"26e8cd8d" , x"7140fd12" , x"1372e9e9" , x"e783d736" , x"973c6f09" , x"087e7216" , x"7bb883c0" , x"884d1a0a" , x"cee62a97" , x"b76c5eb2" , x"f741bd96" , x"2de6b9c9" , x"1a9ddede" , x"5627059a" , x"b2bdf814" , x"300df4bd" , x"7954ff88" , x"5269d1fa" , x"1bb66494" , x"67632757" , x"3807e49c" , x"8c6ed748" , x"6c964cb9" , x"0c7a21e5" , x"306c557f" , x"8d7fda6d" , x"1b9d7095" , x"465a0a5b" , x"62c2517b" , x"3dd30ee8" , x"156680d1" , x"3e3ec330" , x"8dd978fb" , x"2776fe7f" , x"0470523d" , x"f4d7b3c3" , x"ff1c3f94" , x"ef8780f1" , x"ffcb1b3e" , x"d19744f6" , x"a494621d" , x"ba6f5e4e" , x"9a96bc4e" , x"2d01ff42" , x"b992b75e" , x"5c4145bb" , x"c69967f2" , x"30548a3f" , x"3277a968" , x"004e89db" , x"19e28add" , x"5100de96" , x"3a614579" , x"b31a1952" , x"62695467" , x"a010b92d" , x"b43043b9" , x"8b061f78" , x"565f26a5" , x"7064bdf8" , x"f237fdfa" , x"4994d54e" , x"ce878198" , x"806cbb22" , x"89bda905" , x"c2f4b0d8" , x"cec1e63f" , x"c32d2c80" , x"1e099fca" , x"9378665d" , x"4cc39ae8" , x"bf66d4ee" , x"60d888cd" , x"a541bfda" , x"bd08ca94" , x"1f8b5072" , x"cb760515" , x"812037dd" , x"ca2aa1c5" , x"58e61e01" , x"6a718d71" , x"1796fd85" , x"e51ecd29" , x"25d9767d" , x"af7200f9" , x"32bb3fe0" , x"091b38d2" , x"ac19e6f1" , x"dfa16750" , x"6e778443" , x"93600ac7" , x"b1c4747a" , x"127a4362" , x"41bca205" , x"aae746d3" , x"027f8aed" , x"d0e105cf" , x"8843b417" , x"735e20ef" , x"47863b59" , x"cc369500" , x"f23c23ba" , x"5edb6ea8" , x"e80caa60" , x"cab80e9d" , x"6486f9fb" , x"9b9e9703" , x"065ce9bd" , x"03fc3a43" , x"abe3483c" , x"54e0b4cd" , x"d650d08c" , x"a0ed8c22" , x"f8b43355" , x"34fb4cd1" , x"0e93274e" , x"88172718" , x"73486bea" , x"0266d421" , x"951cc618" , x"86c9f18a" , x"afc77ef6" , x"6bab159c" , x"b82cbea5" , x"80918dc6" , x"a6691204" , x"d4b1c5b4" , x"ba17127e" , x"79403d8a" , x"5fb47b0d" , x"53bfcf90" , x"94e2902e" , x"dab5e182" , x"1db9f15b" , x"f6c80dfe" , x"0ec26fba" , x"5f1dff7e" , x"fad1e4c1" , x"55e13bd9" , x"48ea3520" , x"7fedf53e" , x"98503c4c" , x"9ac8301b" , x"f6502f7a" , x"8d6e990c" , x"2f8f2a1c" , x"6d2e1d96" , x"316b0eae" , x"8393d727" , x"5775fce4" , x"8293a1b0" , x"eed26595" , x"085df1a4" , x"6402c9b2" , x"2b0d3a23" , x"45f187b2" , x"cca51e85" , x"26e600f2" , x"d551b577" , x"65a8ecd1" , x"a448c505" , x"5fedcfd6" , x"250e648a" , x"2190bbce" , x"1631d366" , x"6f5ed418" , x"be52153c" , x"176d683b" , x"62a70010" , x"9d58313a" , x"df3e9a59" , x"02cf8692" , x"d2a16315" , x"92c13159" , x"31ab3bc3" , x"ca2bbc66" , x"4729b7da" , x"3c40ff20" , x"89fbf9da" , x"72b16b9b" , x"0a54c41a" , x"91c1752c" , x"c7599d7d" , x"0fb80157" , x"148806f0" , x"7f0cc9c1" , x"a9886000" , x"a46ec563" , x"7221a391" , x"38a4def9" , x"94f8c88c" , x"d64954c2" , x"53b934d7" , x"f89862f7" , x"4802832a" , x"d8abe4d7" , x"06e7f569" , x"81892e31" , x"56bfe594" , x"47646444" , x"ec2a8e0a" , x"bf224e67" , x"330f5d76" , x"3ca77828" , x"d98c4754" , x"f5149481" , x"9c45b92a" , x"9ec95c95" , x"cfc229a1" , x"99aac7ab" , x"5fdb3f81" , x"2c2fcf04" , x"0dc0bf74" , x"1720f6b4" , x"ed00df20" , x"4158dd1b" , x"e212b768" , x"dbcb4754" , x"088a8d60" , x"e93bb0ae" , x"f673f098" , x"b31b32d4" , x"ab4ba05a" , x"b9a58d00" , x"13b1956f" , x"3ad9d077" , x"33fd2ec6" , x"93783d5d" , x"1d2f111d" , x"cf8552d0" , x"81d2070e" , x"67624779" , x"5f540e29" , x"fd0a5b19" , x"b5a4110e" , x"170a298b" , x"78612863" , x"52293111" , x"3955344d" , x"82ebb227" , x"d8e22b66" , x"0f83e610" , x"d2b84bec" , x"b9c6af0f" , x"55da35fd" , x"8e7a7012" , x"13cbe37c" , x"87842166" , x"67c416e3" , x"d479ba9e" , x"4eb26a62" , x"dbd7a1dc" , x"73dd13c9" , x"c9fdcca2" , x"69da1e65" , x"515d81cf" , x"5abc56c9" , x"73c3de2d" , x"075b02cb" , x"c092033e" , x"1401fcaf" , x"1c1fe59d" , x"8a4179fe" , x"1c181365" , x"60c56a0a" , x"4517189a" , x"2aae360c" , x"864ea212" , x"85e6382c" , x"f8ffa93b" , x"b04cdbdd" , x"b5dd57f3" , x"b083443f" , x"4fd60db0" , x"4aba625c" , x"4a9cef35" , x"7b76f635" , x"d9b104a7" , x"cf804835" , x"e961b9b8" , x"fcc5608a" , x"a3a79a19" , x"0d4effba" , x"415ff2a7" , x"30544c0b" , x"16b2cdf6" , x"99b02d0b" , x"d697eb0c" , x"714b0f1b" , x"95b01e92" , x"98c9305c" , x"f2b74112" , x"5c9f66e2" , x"0f9f978a" , x"37ef0e9d" , x"95ab0d7d" , x"6e687a9e" , x"48fcd7e1" , x"7dd50f86" , x"d3e64162" , x"b67554a7" , x"30e47cdf" , x"2632b919" , x"7149a4c8" , x"194ac163" , x"64b69dc7" , x"8dc02d7b" , x"d39a5a2b" , x"7db4c47e" , x"ad476c91" , x"4f67f9f5" , x"352578f1" , x"99b2f455" , x"516f4fbd" , x"9c25b7b0" , x"22416fda" , x"6f99cc0e" , x"abe4fdf0" , x"764953ef" , x"922c789f" , x"db59e8a5" , x"2b75dabf" , x"e42c5235" , x"25ccc4cc" , x"ef7517ac" , x"79e05c42" , x"21fb1f95" , x"e8796662" , x"22870161" , x"8d5b57ac" , x"8b4cab9d" , x"086ebfb7" , x"90c17879" , x"0dc9f5ef" , x"9c0f7f96" , x"ce189fb5" , x"6efb342e" , x"738d4d71" , x"798126b8" , x"61f51a69" , x"8f2e8d53" , x"ca2616e9" , x"d6b75ed4" , x"5d41e77c" , x"f6e9227c" , x"884815c2" , x"c6c8cc53" , x"b62f225a" , x"31595951" , x"df1915d0" , x"40316465" , x"54250088" , x"e55659c4" , x"a66e228b" , x"4cfd07fe" , x"f98edc8c" , x"f50b2e53" , x"137298d9" , x"a292e6b9" , x"9646e353" , x"e5f71f24" , x"69f47724" , x"618a5c33" , x"4f239093" , x"cd663fbf" , x"438aa0b6" , x"9f6ec78e" , x"c23e819e" , x"2e9eced4" , x"fec67973" , x"db454cdb" , x"2fc32563" , x"57a32ac8" , x"c7f922f0" , x"2e416fe7" , x"321fd118" , x"290fa6e1" , x"fe0b3cce" , x"bd9972b0" , x"cd6103a9" , x"27cd4c25" , x"6c9a1f2e" , x"28feba85" , x"ba96d284" , x"6422393d" , x"7f9419ad" , x"9643c590" , x"cf19fc6a" , x"a337b438" , x"5b442b7c" , x"10437218" , x"12c014fe" , x"5e3e583d" , x"974b375a" , x"64f7a765" , x"e90211d0" , x"b18e70b1" , x"319aa4e0" , x"b750b8fe" , x"6eafa7c8" , x"a3df32c4" , x"bfc8ee91" , x"be9e5a0c" , x"0a07fe91" , x"c54b9ba4" , x"f2425ac0" , x"14d1103e" , x"c3801850" , x"6fb53386" , x"8f0edd1a" , x"a62b93a1" , x"2f1054c4" , x"50a592dc" , x"7f7992d4" , x"9cb4e6c8" , x"8491877a" , x"eb0fd8fa" , x"fe86b5af" , x"f7f1348d" , x"dad78f52" , x"ae70a6c9" , x"f6601adf" , x"34d5f4a7" , x"adcf13e4" , x"abc1bdd7" , x"674bddf8" , x"a6714648" , x"ef5aca18" , x"aca12c6a" , x"7abf7fde" , x"536e71cb" , x"3b56b1f9" , x"7ca44a38" , x"6573471f" , x"c895e904" , x"b47ff503" , x"c60ba332" , x"8efdb985" , x"92954ace" , x"c1b28cb7" , x"9bed4bae" , x"fed7d8ac" , x"f2422334" , x"f661e790" , x"732f3214" , x"88fa286d" , x"31ecb769" , x"f6c03144" , x"ee8eea83" , x"1d99a855" , x"cd3cf0a2" , x"0d2bb724" , x"06deb863" , x"4de9d009" , x"00a639cf" , x"948773a6" , x"a608ae75" , x"87ed4949" , x"710d4017" , x"e6b592d6" , x"a6afb271" , x"8a61833c" , x"ef8f8ddd" , x"6e96481e" , x"21159dd2" , x"8aec3949" , x"1d4370c5" , x"b660d107" , x"a06ae123" , x"0444cb55" , x"15fce682" , x"cd0926a6" , x"18f9b729" , x"247b7db9" , x"cf61ba04" , x"7a7d4d84" , x"a8b586b3" , x"41bff62a" , x"b543cbbb" , x"5e7ccaeb" , x"e5d352ae" , x"a9696cec" , x"245b9a6a" , x"2b6b7ba0" , x"97327971" , x"475e63b1" , x"d376beff" , x"32bea9d1" , x"e654ba38" , x"31f0353c" , x"feb11a54" , x"53abc36a" , x"05982375" , x"e15dd27f" , x"7e12ff9d" , x"789a21a8" , x"fa9e336b" , x"676a8967" , x"507a8fce" , x"2de21d2a" , x"8d385164" , x"f80b77ef" , x"95d61b84" , x"684f04f3" , x"63703d90" , x"d8305372" , x"ae3ea8e3" , x"9d85f205" , x"84ae2028" , x"60699573" , x"3bb1fe11" , x"e08efba8" , x"70683f62" , x"c8ec16a7" , x"9aef378f" , x"77073e71" , x"87c4b258" , x"d060caba" , x"c327edeb" , x"e6006f57" , x"d3c5bea1" , x"6de293db" , x"06e30f9e" , x"55969cf1" , x"1af1db8d" , x"98bddd56" , x"c6c37068" , x"e6e8dea0" , x"057f8af8" , x"b3baa06b" , x"bcf2fdaa" , x"60a0e5d7" , x"38d257eb" , x"bc261253" , x"7dc95f88" , x"f4401490" , x"4754a6e2" , x"8af5ccc3" , x"c4f5262b" , x"8a44602c" , x"b2e60fe3" , x"4fa4e189" , x"fc8e6851" , x"123c6dd6" , x"6615ce11" , x"2e96459a" , x"d8039532" , x"17ce1f4b" , x"7e65c7de" , x"76a73b3a" , x"c97de704" , x"02639d86" , x"8f9722ae" , x"ea3f2357" , x"ef2eb1cb" , x"a48ab8e1" , x"eace87d8" , x"005cffc3" , x"c490439f" , x"07c7544a" , x"3d2a6f7b" , x"355e4de7" , x"ba4a1126" , x"7478a94a" , x"4c91d22f" , x"209481b3" , x"d82f4c38" , x"0236bc25" , x"04fab43f" , x"ba21e394" , x"242c5622" , x"5aa76077" , x"85814bd7" , x"c7cb4e33" , x"b639c3b2" , x"6fc8bac1" , x"5b3cf6cb" , x"6fc20df6" , x"099c3da7" , x"0c993c28" , x"414e5aae" , x"0cb4ad23" , x"0ee99fa2" , x"17525749" , x"9078b040" , x"9812cf8a" , x"b552ca2c" , x"3db7af4c" , x"244dd81a" , x"d763f72c" , x"46ae9580" , x"db724bbe" , x"9bdd020e" , x"f6af4a04" , x"48e6b489" , x"7d288958" , x"84a645b8" , x"38663e32" , x"275db211" , x"39e8cf38" , x"d3e330c6" , x"896aece9" , x"8a319eba" , x"c3199f26" , x"a8352468" , x"58fa293e" , x"42bb0cd7" , x"761348da" , x"d3b4490e" , x"a3aab8d1" , x"d19d869b" , x"ead688f9" , x"37b8c511" , x"295cd1f1" , x"c650ed2d" , x"b733e1d3" , x"0612842c" , x"93e6b1e2" , x"56fe57cb" , x"6eecae9a" , x"4406fe84" , x"e25dbc30" , x"48ff2646" , x"649f0a2e" , x"97d5781b" , x"2dd150cd" , x"5aa96822" , x"a2222658" , x"3777d4fa" , x"9fbe801a" , x"aba8bbff" , x"53f3fb1d" , x"0ffc245b" , x"cd8f2283" , x"5ee74a51" , x"ffddc7e0" , x"5f56908c" , x"fb21627e" , x"fa59b049" , x"20857e33" , x"c0e2d2cb" , x"3b74170d" , x"bdcb17ab" , x"060cc6fd" , x"fb5dfa30" , x"9b80b416" , x"e1995975" , x"1c5dfff0" , x"58298154" , x"684f4438" , x"66417da1" , x"e252db96" , x"5e1f3663" , x"8c526e04" , x"09054d59" , x"5e76fc59" , x"94cc5713" , x"35562995" , x"737d8c41" , x"70e1a889" , x"c08122a2" , x"f4c94575" , x"114060c5" , x"1fc02995" , x"bee0cde1" , x"7883f0b7" , x"4942540a" , x"db5d8ed6" , x"3f189c03" , x"0b1ba348" , x"82b46479" , x"b10e586f" , x"9dd8cc88" , x"fa9ecaa7" , x"1507595e" , x"48843eb1" , x"c03e35bf" , x"223f705c" , x"c28c7150" , x"af6e7d5c" , x"495356f2" , x"e8d20382" , x"31228736" , x"9c61e8dd" , x"ebd08c5a" , x"e66545d8" , x"2d2254a6" , x"3184dfc7" , x"b42af5dc" , x"c121f838" , x"4652fcca" , x"58a48ad3" , x"afb7c4d7" , x"6b2b08fa" , x"fda306e5" , x"27dd413a" , x"d5b414ec" , x"d1aa05b5" , x"9af729d8" , x"9ffafd0d" , x"14ce3f1e" , x"bd124bb6" , x"c7806ae7" , x"ce1bd8e7" , x"e4516e28" , x"11358111" , x"5e45c0e9" , x"f366fe98" , x"15f58bec" , x"7f6134ee" , x"eca72421" , x"c1513dfc" , x"a32d358b" , x"be0e4227" , x"d7894910" , x"d4c4e862" , x"534e6c26" , x"28108149" , x"4c721d25" , x"75122f25" , x"778d1d08" , x"9e3bd58b" , x"42ef1669" , x"eea3916b" , x"fe6bcdfd" , x"d5c857ad" , x"a80399ea" , x"e53a79bd" , x"f613e5cd" , x"951fef0d" , x"e61b5bf3" , x"952ee510" , x"5960f344" , x"dadc6d28" , x"23063e60" , x"08ecf574" , x"0baa0076" , x"e2aae429" , x"8aa09e9f" , x"68610be7" , x"22c38ef9" , x"0950553c" , x"777bef48" , x"bf038d3c" , x"a04a1df3" , x"27a2dbb8" , x"d6d8d7ff" , x"24d72d14" , x"ea3e9f2a" , x"9b2021eb" , x"65ecc71b" , x"4125a815" , x"b545d858" , x"52fbc519" , x"eae317e0" , x"66dbc50f" , x"1fdc8861" , x"680814fb" , x"eb13f1be" , x"62dd6c3d" , x"30fe3456" , x"9c1bf8ec" , x"5366bf1d" , x"2ab959bb" , x"9edbd0e4" , x"3026cd42" , x"b8155c4f" , x"183998f6" , x"ea8605fe" , x"52bc55f3" , x"4034c52e" , x"c5044df4" , x"529d170d" , x"3bef2843" , x"5fbadf4f" , x"bd889775" , x"38fdb93c" , x"b15c8c35" , x"6bca7d0b" , x"d2f6ca20" , x"7e09a776" , x"d3f6562c" , x"7b02b91e" , x"4b1a292f" , x"9216cb4e" , x"4f32d29a" , x"d4c08497" , x"85e547f4" , x"392278df" , x"5346cb78" , x"b17b83b3" , x"d4f3a162" , x"cfae7d02" , x"cf6f7aa3" , x"d2e96342" , x"8e97703a" , x"20f6c2dc" , x"43519c69" , x"27298162" , x"ae399631" , x"6d48c5c2" , x"3bd0b153" , x"5242b6b1" , x"74d84afc" , x"70a022c9" , x"6272f9c9" , x"d8690408" , x"89e1c8a5" , x"664adc1d" , x"fde04b98" , x"46d32915" , x"c1561fc7" , x"73d37c5b" , x"faff16d7" , x"4c1082c4" , x"3c1ab71a" , x"9a860b34" , x"874fa5ed" , x"fab2b7f0" , x"0d2ae9db" , x"3f3dcb89" , x"c1c29754" , x"18303ad9" , x"9a1b5897" , x"880e6b3f" , x"db6f6887" , x"a6ace660" , x"fcffbb13" , x"43fbfbaf" , x"edf2b1de" , x"19a9a890" , x"68d5f871" , x"f2bf230f" , x"001660ce" , x"487a51ce" , x"8a77007c" , x"9b0f9246" , x"352dd587" , x"1ece7750" , x"3822f801" , x"fe583563" , x"53680a0b" , x"5a3427e2" , x"1890240e" , x"b332e717" , x"bf5e5dae" , x"ae99e23a" , x"bf9e4863" , x"a623520f" , x"8b15abe0" , x"88497d1a" , x"568fd6e6" , x"4988404a" , x"d513d1b8" , x"002929ca" , x"8d755ecd" , x"4a6866cb" , x"f5218bae" , x"9ee4ee3c" , x"e490b97d" , x"99ffe192" , x"5b43d234" , x"83bac1be" , x"8be0fe8e" , x"a6fb2eb9" , x"58c02287" , x"fe1481e1" , x"9f7000e3" , x"8de8726c" , x"cbef9865" , x"54afd3d6" , x"bef1a852" , x"a831ca73" , x"2023247c" , x"c10e6b70" , x"d28869e3" , x"1ba6b2ec" , x"06704364" , x"28e847f4" , x"6a1802d1" , x"d0b1585b" , x"bb3d8519" , x"97f39335" , x"c808207c" , x"090a2606" , x"5e067328" , x"0e2a5083" , x"beafa8f4" , x"533268ed" , x"e46b9f55" , x"c5f8cbd2" , x"3e1b417c" , x"4fc2a2ac" , x"212d4476" , x"a70fd8c9" , x"399e0c6d" , x"c8f47898" , x"599a8302" , x"fa0650e4" , x"497e609c" , x"852e5cee" , x"ed6fdaa7" , x"122491e9" , x"0d22e5e5" , x"dae77e5b" , x"97b90229" , x"584d8dec" , x"29b3be0c" , x"47ea8da8" , x"d6a1c2a5" , x"8c2fde93" , x"2ae545f3" , x"5ac20a8e" , x"80903834" , x"99b7d39d" , x"ffd40e81" , x"32c0e2ff" , x"5afbf69a" , x"5bae3bda" , x"0c0d48f2" , x"3710089b" , x"36b275d1" , x"4c4df09a" , x"65d8c8ea" , x"58b92602" , x"556b4735" , x"1397f392" , x"3ac73b44" , x"2f0ec08d" , x"efa59262" , x"5bfa0ef0" , x"aee575cc" , x"7a3e4833" , x"f64d16fd" , x"bd47ee85" , x"701f0283" , x"d3aa1ee6" , x"f0b9e73a" , x"4fbe282b" , x"017e5ba2" , x"c9dc5417" , x"9c3d14ca" , x"f55a1e46" , x"cd134d01" , x"0e4dad26" , x"3ba4ad86" , x"14ab1c54" , x"eeb64477" , x"1d000d91" , x"c3653077" , x"92803d5d" , x"d3923263" , x"8689c580" , x"92ce827e" , x"f4099f6e" , x"cae6a1dd" , x"3671ec91" , x"543c0b39" , x"b95494d7" , x"3934cdd0" , x"bae16c27" , x"4ff88d33" , x"1584a36d" , x"95a354b8" , x"4031c6bf" , x"d47540d6" , x"716729f9" , x"4a5bbff5" , x"af481352" , x"670dcde5" , x"e62d9d96" , x"dcafc989" , x"006346c3" , x"9d5f9223" , x"bde5c1d8" , x"fdbe7b8b" , x"f891788f" , x"34259c00" , x"393bdea5" , x"d3c3f978" , x"f6665635" , x"ad054457" , x"f030b354" , x"3fbb2714" , x"416b8906" , x"79cd1628" , x"d02f20a5" , x"6629cb59" , x"3b7b9c1e" , x"9974c8f3" , x"de8d8d37" , x"ccef0f59" , x"d6a5e703" , x"1ae5c976" , x"c4363c7c" , x"d24a0914" , x"fa9e62b5" , x"d7516f0c" , x"454313a3" , x"5ac0ebcb" , x"af6bddc4" , x"6e19084c" , x"278be084" , x"927e44f7" , x"c4919342" , x"b3693ffe" , x"171fad0a" , x"be127f63" , x"e43c48fa" , x"c204b216" , x"c895871a" , x"639df15f" , x"8bb3b42c" , x"6de6c493" , x"2953a037" , x"f4d300fa" , x"1d5b71bb" , x"92ae406a" , x"1fc4e267" , x"d9876261" , x"8c791fa5" , x"46be910b" , x"7f3aaaa0" , x"9f5099a5" , x"b4ddb9fb" , x"969edf1a" , x"8d13b1ba" , x"f6a5de8b" , x"7af2537a" , x"15fdb812" , x"8c2e4c99" , x"8020b21c" , x"18fc590f" , x"8586e6a6" , x"53ec44ef" , x"17151e70" , x"f436cfe8" , x"e79838f5" , x"8073c921" , x"e2675023" , x"fec08616" , x"7061a069" , x"b1b21143" , x"c81ef931" , x"082ee456" , x"2601cddc" , x"11227752" , x"9eac41be" , x"8900bab8" , x"42b83bd8" , x"1c7f7069" , x"72168698" , x"2b234d25" , x"d8105a0e" , x"dcffa585" , x"323a7c5e" , x"6a1eda8d" , x"4dc93858" , x"7555161f" , x"7bb9315f" , x"d60694d7" , x"567ad9bb" , x"04f7bc38" , x"cc69913c" , x"e0ea773a" , x"fccbfc4a" , x"c5282a47" , x"28b7573e" , x"7054e664" , x"3ca4274f" , x"5050d80d" , x"b3c5c7ba" , x"5ae4df99" , x"601ee92d" , x"7ee2bb8b" , x"f944b975" , x"c78d25bf" , x"f8e90441" , x"9b354f0b" , x"a4c96521" , x"b61c84eb" , x"dc2f70a8" , x"1b51d239" , x"66e1d484" , x"9a0029b4" , x"a1c6376b" , x"f52fd80f" , x"fc3877e8" , x"48dc72e3" , x"8f39e95d" , x"4c87b4d8" , x"eeffe12d" , x"d2d17421" , x"b8686989" , x"7d5a1ed2" , x"7be9f2a7" , x"fdb4f329" , x"a3978abf" , x"618b52c1" , x"e33c2b7f" , x"6dc2202f" , x"32e06977" , x"11816a9b" , x"6536b96c" , x"04a1cd0b" , x"fdff3346" , x"e0ee1118" , x"670083e0" , x"e1dc665b" , x"a8aad172" , x"f7ba20af" , x"e6bec034" , x"35f42574" , x"fed15708" , x"896dfb8d" , x"a735b56c" , x"99ff7d24" , x"1bc27d59" , x"faad0e16" , x"093ec4f5" , x"298ad608" , x"9e3b3a25" , x"cd34fba7" , x"91305f7c" , x"b3b39177" , x"f64350cd" , x"c97422a7" , x"bf00c48a" , x"f42ab3c9" , x"a99aa7b0" , x"7ed14aab" , x"85f7dc97" , x"a1206432" , x"42886e63" , x"fb24abac" , x"f6453936" , x"bee2effb" , x"8a4acfd9" , x"924d4348" , x"07bfc90c" , x"8f75b955" , x"b241aa38" , x"40a91ff5" , x"850c1e24" , x"ebc89647" , x"0f1ca065" , x"10596e2d" , x"e3d96a38" , x"0fc2fa71" , x"54882247" , x"c54f028b" , x"3acdb28c" , x"e5aaf94e" , x"1d2bbcf6" , x"d657f616" , x"4f98a187" , x"2eef3d54" , x"3a7a8a6d" , x"4760ee24" , x"a6e9495d" , x"7240dd41" , x"10efdead" , x"9b97c136" , x"4682abc8" , x"065bbbb2" , x"48255ef4" , x"fd662448" , x"e14c05b0" , x"deb10eb6" , x"71bfa266" , x"39dd8427" , x"c183967f" , x"df130322" , x"9a71a18f" , x"df60c30d" , x"c8841ddc" , x"89c4da33" , x"1d2a8efe" , x"791700e3" , x"fa8329be" , x"5e786ef0" , x"d93da1be" , x"c56e916b" , x"0cf72b21" , x"d9372423" , x"775900c7" , x"ebba6310" , x"535e0344" , x"ade594ff" , x"a1551f80" , x"0d2a04ce" , x"3af4e2ce" , x"85c5227d" , x"94735768" , x"9d7ad19b" , x"9a6873c8" , x"f55206d2" , x"9991ad2e" , x"513fd6b4" , x"72cc2b6a" , x"46e87b04" , x"09118305" , x"692655e3" , x"83895e77" , x"c58323a7" , x"686100ff" , x"f340081f" , x"1ba8e7a0" , x"8dcf5922" , x"75ba68c3" , x"144700f2" , x"736d0d43" , x"caf1e69d" , x"8d178877" , x"ae4a9f70" , x"ce2efa3e" , x"8cda3f8f" , x"b36ae916" , x"701f6fec" , x"df4ad370" , x"9e06d89b" , x"0d5c770c" , x"1e51df7a" , x"383d08cb" , x"803a114f" , x"75ab194b" , x"4a5e401c" , x"f5627534" , x"7bee52b1" , x"ca40698a" , x"d4aaaa6d" , x"73ae0df5" , x"5dd7b5c5" , x"555b8cac" , x"a34fe55b" , x"0f20decb" , x"9a767510" , x"bdabf849" , x"6ae330cf" , x"81bd4932" , x"94e1d49f" , x"332e4fdb" , x"b895213b" , x"6d5c8e71" , x"d8564c0e" , x"2b2f4921" , x"f1c754fc" , x"c06f0e9e" , x"226869a2" , x"5e4c3db9" , x"11ff8966" , x"f11af890" , x"aac4deb6" , x"04656b64" , x"6cce57a1" , x"d43d021b" , x"76158551" , x"a0684435" , x"0b369c5b" , x"89eb4aa6" , x"3b794ac2" , x"a687ab1a" , x"de0b93be" , x"ba046494" , x"ec839792" , x"1830671d" , x"5f144140" , x"e0a8af76" , x"9d633a9b" , x"03ad3cc4" , x"54633b9d" , x"4b576aa7" , x"eb73ac1c" , x"2e0ee6c1" , x"39ea8c27" , x"ed219f0b" , x"230f413d" , x"117445ee" , x"53315f7a" , x"94c28684" , x"c3037eaa" , x"a31c57b2" , x"7ad16d35" , x"a6b9952c" , x"0871719c" , x"dd57de5c" , x"19ddd2fd" , x"0e52e7ae" , x"5f73fc3b" , x"d11d6ba6" , x"876aaaf5" , x"8767767b" , x"b8008976" , x"b1c0f55e" , x"aea945af" , x"36602adf" , x"98537472" , x"8b146513" , x"0db9da6d" , x"b3d85e47" , x"cd68bf90" , x"f4d8e53c" , x"4195688b" , x"71cd83fc" , x"19e09811" , x"15dca1c7" , x"d3eace4b" , x"0eadd810" , x"5380086a" , x"a123aad2" , x"21fd1059" , x"cbd2642b" , x"62f72ad6" , x"b0f1ea57" , x"4f3c29d4" , x"58661899" , x"ba206103" , x"f26293ae" , x"e622563c" , x"852b315f" , x"a3502268" , x"f42d1734" , x"2dca9696" , x"12d729ee" , x"07657833" , x"35000ba0" , x"b19bb226" , x"c6683912" , x"5457e774" , x"ea08368c" , x"5525e408" , x"c8553d3e" , x"fb08eae0" , x"4ba82104" , x"5b05b77c" , x"26df5c72" , x"db06924b" , x"d910a9fc" , x"da2d0030" , x"c8ec3b08" , x"06e25de2" , x"45553696" , x"e3bb5076" , x"3a51cd7a" , x"36e97b18" , x"522e93df" , x"d53ae31c" , x"d45e298e" , x"9f3dcb82" , x"d27a8848" , x"29514ddd" , x"92184579" , x"99a96bdb" , x"92636d51" , x"93e44e17" , x"49387e4a" , x"b38bc93b" , x"b2fa6ab1" , x"e5e0cef5" , x"cbd78f88" , x"0c98c62f" , x"710bfafc" , x"d3873030" , x"723b2fa9" , x"996d6ded" , x"7735a6dd" , x"773cec1b" , x"476f1caa" , x"bd2cd4cb" , x"ace56582" , x"c8ffb708" , x"e7568ef2" , x"9a4b3b28" , x"e895272e" , x"f8fb7097" , x"bf484c97" , x"35b34e53" , x"42b0e1d8" , x"993e786c" , x"b08c1b05" , x"099e77ae" , x"21bfa798" , x"669e3103" , x"1f9dc035" , x"1ebd1429" , x"30df0260" , x"3b2f77af" , x"254eb2e2" , x"4a830d1a" , x"95c56b07" , x"d2807db4" , x"12c7d4fa" , x"5d662e0a" , x"d283f8a9" , x"376ed66b" , x"b9102b42" , x"a2f429e8" , x"ed050848" , x"5030cbd8" , x"7e1d9020" , x"692000a3" , x"a7a667c9" , x"bc687ae9" , x"e3df21cf" , x"d9fa4fab" , x"89dccff7" , x"133b832d" , x"483e990d" , x"0451a3ce" , x"f9d85a1c" , x"aca3647b" , x"09532eb1" , x"ef60015d" , x"5384c3a9" , x"5e550ae0" , x"f9176bbe" , x"e974f534" , x"5d72c724" , x"9d4a272e" , x"4f246df5" , x"75d4a41f" , x"1ef41d2c" , x"8ba431ed" , x"ea6f9f1c" , x"2d3a9617" , x"22aeb300" , x"f5c851ce" , x"5505ad86" , x"de8db308" , x"e5c13e1a" , x"15669be2" , x"7fe8fb73" , x"c2b92839" , x"9d8387bf" , x"ef6a7c90" , x"954833dd" , x"1947ffc8" , x"b2c0c4fa" , x"9958bb89" , x"07825302" , x"66c2a854" , x"872351cd" , x"ffb25218" , x"0835ed17" , x"93b52efa" , x"d3bf9967" , x"4dc16c9a" , x"5709560f" , x"2f74c5a8" , x"d8c20cb2" , x"2c741386" , x"3efe6a5f" , x"3a17b23c" , x"94dc9c41" , x"bea652ae" , x"f00b9798" , x"4ebb6811" , x"0c3bc9a1" , x"cfaa7e8d" , x"0dd17ac6" , x"c6ce752f" , x"05473921" , x"b2067f8f" , x"ae75602a" , x"db31fac7" , x"993fb806" , x"c2bd4067" , x"1d31128f" , x"280d4c6f" , x"cbd6bc25" , x"e7ad2b46" , x"9e2b74db" , x"0c9eed1f" , x"11f98377" , x"aa1651ab" , x"11bc4443" , x"4bd722e8" , x"22d1614d" , x"b119e711" , x"c9f4c812" , x"903379cb" , x"17a76cf9" , x"17de93c6" , x"3ce4f812" , x"d348838f" , x"3e5fb5a9" , x"436c0bbc" , x"1ad5a0ea" , x"3a1d4eee" , x"dbbd01a8" , x"4ce92770" , x"b2bd385f" , x"4e875736" , x"bbd6864e" , x"1081290b" , x"a6892cd7" , x"68a47875" , x"842a4ed6" , x"5f193154" , x"538e2c28" , x"f012cc3a" , x"a96a2a29" , x"937ab976" , x"1e18c583" , x"3cb5eef5" , x"25d75cae" , x"7d83a86b" , x"050f4c0b" , x"42a755c8" , x"f6dbd2ba" , x"2b84d545" , x"f86a5bca" , x"389305ca" , x"1fb55278" , x"dbb1492b" , x"77a82eea" , x"d68ce11c" , x"a81d192d" , x"1d60517f" , x"4a4999f6" , x"73acd677" , x"c129503d" , x"79b8c5c1" , x"8ee0d305" , x"cf26f9e1" , x"6d83d0d3" , x"3ad00613" , x"4466d46b" , x"4d6d0972" , x"c0f4d8ec" , x"61bc45d0" , x"e5fbfdbe" , x"3b32e5f3" , x"ba7b4ee3" , x"3685213f" , x"6826051c" , x"5af24967" , x"f035779a" , x"39aac846" , x"4163b19d" , x"abaac0da" , x"887d62dc" , x"cec111c1" , x"f46ad0b7" , x"7fb4b1a5" , x"448b1a5b" , x"04c21ceb" , x"40058bab" , x"95519f9c" , x"ed7bf588" , x"d68e0a0b" , x"118e9ce7" , x"010747ed" , x"4ca580ee" , x"a58266db" , x"977204aa" , x"e06df822" , x"340b69a9" , x"64e1b851" , x"a2c93ddf" , x"3a5c40ba" , x"cc61fe47" , x"1bd7238e" , x"806f7ae8" , x"622f4f91" , x"a69b9fdc" , x"3dee882a" , x"cbc3b4b0" , x"c069eae7" , x"3bbe6201" , x"ece4b3ba" , x"99d094b7" , x"35ed23f8" , x"1cca5597" , x"e97e2445" , x"840937de" , x"27032279" , x"d67cba20" , x"f45d9913" , x"ebb8e699" , x"42ad8eb0" , x"7f8bdd84" , x"b7b76567" , x"471185db" , x"190d1e6a" , x"a70b8c49" , x"9b358211" , x"ead41825" , x"57decc25" , x"8284d6a0" , x"18734e03" , x"f9649ce6" , x"97ca7d71" , x"3280df73" , x"63fac25e" , x"1c769e79" , x"e9702614" , x"4c1f6920" , x"aabf53b3" , x"657baf71" , x"2e206b0e" , x"6bb6a4f1" , x"dcb407e5" , x"4fbcd94f" , x"d4f2e30a" , x"b19fb4a1" , x"fda7a0b2" , x"1784e986" , x"ba98e4f5" , x"66ef4781" , x"e6dd03cc" , x"4b90f802" , x"ddb9b2a7" , x"4e7692b3" , x"51fb297e" , x"1b060de7" , x"21e4f028" , x"980515ed" , x"e8864060" , x"4860d48b" , x"df9ab7ca" , x"27bc9aaf" , x"4c89c110" , x"002b2a99" , x"ddee285e" , x"4899b588" , x"8d2d5191" , x"8d01f118" , x"328c5758" , x"def37220" , x"742f3580" , x"0ad11edb" , x"bf9386ef" , x"e79bdc13" , x"d2f62763" , x"21878492" , x"4c7eb549" , x"d56f42b0" , x"2f561d1e" , x"cceb7ec0" , x"9d63d230" , x"eafa3080" , x"8644de6a" , x"2326553d" , x"152b6929" , x"81362306" , x"e925f244" , x"67ab5be6" , x"22bbb768" , x"2c6f39a9" , x"2a4d1605" , x"933f3bbc" , x"a5f4e069" , x"9b311939" , x"9530d181" , x"36e5ea8a" , x"0ed336fd" , x"851a47be" , x"fcd2ce6e" , x"fd3b47eb" , x"f08c2dfc" , x"7d6b1487" , x"030a5bd9" , x"b1e335fb" , x"a751f6af" , x"6952f0dc" , x"ebed954b" , x"08e720fa" , x"0b1e85ec" , x"4af70244" , x"20f92427" , x"cd2b4921" , x"2b3b3a34" , x"58b45ab5" , x"ebbd116c" , x"15543196" , x"d207edcf" , x"82d7ddf3" , x"dfd08b35" , x"5de8cb46" , x"8e7247ff" , x"bd4e8771" , x"0c6ea650" , x"86555f01" , x"983a76ba" , x"cdf51491" , x"4d13672c" , x"d1211754" , x"6e094b07" , x"308133e8" , x"cae8b344" , x"1faa5fd0" , x"bfb1695f" , x"d22cd346" , x"1b2e4324" , x"a34d422f" , x"4129ae8f" , x"04206d7c" , x"2f378747" , x"e55d4841" , x"834cd36e" , x"83ef9eb6" , x"3c0918ae" , x"8b65ca3b" , x"693698a5" , x"9b3fcbe7" , x"5abb475f" , x"c2abf2be" , x"728a3ebf" , x"daf8032d" , x"cb93d83c" , x"6203aab7" , x"420a9e7c" , x"15ab91b1" , x"c5f38ba3" , x"bbdf1edd" , x"cd62b65f" , x"54fd40b7" , x"f1f13eab" , x"d6f9d342" , x"a8f1472a" , x"5f294239" , x"d8bc83cb" , x"d405ea7b" , x"d6bcec1d" , x"2d30532a" , x"543280de" , x"212836a5" , x"7a9c61c1" , x"e1400ce0" , x"562d47d7" , x"0b48c51c" , x"79a3b756" , x"afcce218" , x"a71189c8" , x"bbd88a9a" , x"2b0ba9d9" , x"6fea887c" , x"456d67d2" , x"613d1f85" , x"6eee3bba" , x"facad46b" , x"cb649b4d" , x"66246eca" , x"ab7d0aa9" , x"70b016fe" , x"87500e61" , x"28248fd1" , x"66106f54" , x"5376fb8f" , x"db853630" , x"50665cd9" , x"8491d9fc" , x"e4fdfed7" , x"cdc0a53e" , x"3f3cfa12" , x"1a15143d" , x"4f88a8e6" , x"a72fb3d1" , x"68aba1f4" , x"e3238b99" , x"b54033aa" , x"99bc1082" , x"24c56ee7" , x"aa0d8a40" , x"df0ef689" , x"21b6cfdb" , x"1549b478" , x"88348ed6" , x"76347368" , x"98ef5371" , x"07c79339" , x"b6419152" , x"c0d1c003" , x"3a83b39c" , x"b335ff17" , x"9b7958d6" , x"36ea465a" , x"4eed3f06" , x"ae0e3bd1" , x"25c31147" , x"8eaabba6" , x"6ee84636" , x"d9c617a9" , x"902c5d22" , x"8efe25ff" , x"3fbd8aff" , x"e6daa389" , x"5bd3b5dc" , x"6b658323" , x"16a3196a" , x"5bae4cb5" , x"d7fe7cc1" , x"7d2e4932" , x"9a60835e" , x"4186bc26" , x"04f2ca9b" , x"edde0997" , x"362a20be" , x"777d5ffd" , x"21c0730f" , x"4106a888" , x"988dfef0" , x"6e645517" , x"43ee08fc" , x"b3d901a3" , x"f64c70ea" , x"66ff1713" , x"c9a6cf8e" , x"2e8d1256" , x"37c503ae" , x"db3345ef" , x"681ba46e" , x"958e3634" , x"0d57be75" , x"5fa2dbf5" , x"70b79b5f" , x"38c0f944" , x"609311fb" , x"380fff8a" , x"ecb5a892" , x"85b10671" , x"fda33ce9" , x"6ef4ca63" , x"de302802" , x"bdc61938" , x"1117dd29" , x"1208fca7" , x"96ed0f14" , x"d8ead81c" , x"b110c6c1" , x"ae0ca194" , x"64fbf26e" , x"22fb981d" , x"cc0633aa" , x"dbc03ef3" , x"76150fef" , x"33285440" , x"308f1a16" , x"9b7aa10b" , x"6c4289d8" , x"8b04fef4" , x"e86b6bed" , x"298e1c76" , x"5ce72a38" , x"01727aa3" , x"f5d09ccc" , x"c5800ce5" , x"a366c480" , x"c3c91e0c" , x"34091aa7" , x"6bcb3372" , x"cdeffdd8" , x"0e8b4f1b" , x"121b9bd1" , x"95f383df" , x"e217182d" , x"2c957023" , x"3a2b1ca4" , x"ba863a65" , x"7531aea1" , x"88c74c5d" , x"d0567908" , x"40c8d23e" , x"bd6c3d38" , x"eac43b3c" , x"33b3974c" , x"c219096a" , x"29120c46" , x"e3147238" , x"8bbae118" , x"119cc1d1" , x"3752130a" , x"2efbb436" , x"6d7cdbf1" , x"bcb0cb29" , x"11cd6bf6" , x"b25be780" , x"9624e470" , x"c6e901c4" , x"79d9eb1d" , x"807cbe19" , x"9820951c" , x"6ced5c35" , x"86958ac0" , x"9c7a095a" , x"f6364562" , x"db13ddc2" , x"f1e0b624" , x"abb95bf7" , x"ea923d89" , x"860a20d8" , x"a3d775aa" , x"4c7f2aad" , x"6f9a999c" , x"b4375146" , x"519df7f6" , x"61b1401b" , x"c15c7d94" , x"9153cdd1" , x"9fe5d231" , x"e34adb0a" , x"33a804f3" , x"d7cb8640" , x"635ea76b" , x"e617a98d" , x"17ee2706" , x"f06281bb" , x"84d8c899" , x"d0c05bbe" , x"f61fe8c7" , x"0058fc91" , x"b1d62960" , x"00ca8d44" , x"6772f991" , x"16645b27" , x"cc1229db" , x"42bf0713" , x"b4c31769" , x"05d6223c" , x"c65c5578" , x"6c90d28a" , x"dc02bdad" , x"575008bd" , x"3a360e7c" , x"8a962bd8" , x"f8f0c12d" , x"ed196ac6" , x"0215c090" , x"4c6a75ae" , x"97f2b94a" , x"568cb98e" , x"e6ede417" , x"dc06e363" , x"402039fa" , x"57299622" , x"4de0fd1e" , x"235bdbc3" , x"b0156c3b" , x"81ff1ccd" , x"11758a9d" , x"db4dd6d6" , x"01404879" , x"62626088" , x"a1b4c53a" , x"b218ccea" , x"96d3f46c" , x"a0be5405" , x"250eb289" , x"734ca35e" , x"cb941c92" , x"793f068d" , x"20e88292" , x"f31ff4bc" , x"08cf06c0" , x"156018af" , x"097283d2" , x"47a2de2a" , x"df01dee5" , x"726f1229" , x"7552f763" , x"966b120b" , x"176f1ca7" , x"e0aca19d" , x"12bf8141" , x"7816f8c0" , x"075c9e6a" , x"6ffaa82e" , x"fe70c3ef" , x"bf05f9fc" , x"4fad6ea4" , x"77c8fae2" , x"a0cd9c43" , x"dc5f2e6f" , x"425df870" , x"776d54da" , x"62f5034b" , x"7f83c68f" , x"91768ed6" , x"7cc84146" , x"fe41fabf" , x"3abe772e" , x"97f7a697" , x"15e6c04c" , x"425fa005" , x"11400862" , x"41f88eba" , x"e36d9698" , x"d8636423" , x"3bb0e0a2" , x"037b48b9" , x"dc918a27" , x"5c0a7dd5" , x"b6344560" , x"1f1384bd" , x"df70ac13" , x"e524b9e9" , x"f020e656" , x"3a6adcb0" , x"23c2ad24" , x"97b4f060" , x"64d6a3d8" , x"8032a1c5" , x"fb062a6d" , x"2a651e0b" , x"a51138ab" , x"321b5ef4" , x"e57b1c63" , x"f48dc28d" , x"7b7373ab" , x"63e728b9" , x"039b9a92" , x"884b9ee9" , x"9f75160e" , x"a5596b8c" , x"3b2910c2" , x"968e7a1d" , x"8705e992" , x"27671084" , x"b99912b2" , x"df234d3c" , x"9b7f99f3" , x"7054eb08" , x"969f2efc" , x"9608ed3b" , x"6ef595f9" , x"771c9f79" , x"3e821d75" , x"01757b1d" , x"6dd05896" , x"160e9b45" , x"029afd4c" , x"f4faef97" , x"9bdbb8e6" , x"a5fda8e1" , x"f53ddcaa" , x"3d7f2d0e" , x"186f2ef7" , x"894ca74d" , x"091c7692" , x"8e1c91a5" , x"e2e04def" , x"1db02c26" , x"3f378c8a" , x"f79cc39b" , x"024841cf" , x"986691da" , x"d09e9d74" , x"55bbf22f" , x"23f7c56b" , x"28aac31e" , x"e13eed54" , x"8ef11b89" , x"186a9ceb" , x"88737d74" , x"5a4160fd" , x"c5e61af0" , x"97ea6913" , x"5b5e430e" , x"95ce76af" , x"fbe1cafe" , x"aaed313f" , x"6a76d626" , x"a5e51ae1" , x"10af10aa" , x"6ef14673" , x"9a89c733" , x"23c73af2" , x"1d496da3" , x"c07e73d4" , x"2d33edff" , x"3de5bd4b" , x"187e9468" , x"a6848094" , x"6b5f6da2" , x"db7cddd3" , x"7dc830b7" , x"15994d80" , x"ef18a30b" , x"f8dad5c3" , x"b2d259d3" , x"080dc227" , x"12e2a70b" , x"d5dd1291" , x"b8b8d510" , x"d5f14f55" , x"d9cbcaad" , x"0cc37618" , x"8deab272" , x"8bbf32df" , x"b4303521" , x"f1739409" , x"ff269865" , x"524c0f25" , x"0d173208" , x"ce749bca" , x"1cd0ee0d" , x"99f544d5" , x"8d53cff4" , x"ca249119" , x"cfa564dd" , x"cc9763e0" , x"a7be5c54" , x"0cb046c3" , x"3989e0b5" , x"487fb4be" , x"34f32e17" , x"a748f257" , x"42bc5e36" , x"7d5a0d78" , x"f3fa9d1f" , x"f90cd81b" , x"ee6a2af4" , x"bf9d08e4" , x"25e6814e" , x"915e0980" , x"fb9c1763" , x"4c88ea5a" , x"c5cc1a9a" , x"41906915" , x"eec540ed" , x"e2f5d847" , x"3685a806" , x"72618a96" , x"abd04e7a" , x"d0e48a67" , x"36e17136" , x"192ca226" , x"37c2c54c" , x"dc0e5116" , x"5441854f" , x"0712b1c1" , x"b3c90a7c" , x"e62f1da4" , x"b8f3d577" , x"e6622c40" , x"3a278e8d" , x"862bcfa0" , x"d78c90e4" , x"1ec5653b" , x"7e8443c2" , x"2d83e9fe" , x"0e63c194" , x"b4c377a1" , x"0ef94cb0" , x"d4d3fe33" , x"a724aad7" , x"08eade88" , x"4110a5ba" , x"c201b7be" , x"e600cf99" , x"f5054dad" , x"f8f25769" , x"57c65cb6" , x"8564a2b9" , x"a363f092" , x"96dace7c" , x"57cf3a8a" , x"c600f767" , x"376aab5b" , x"f8fcdf1f" , x"c94471b5" , x"e986ed62" , x"b91c6c70" , x"8282965d" , x"4761fc9e" , x"475112f0" , x"951a39eb" , x"13961d1c" , x"6bc708f5" , x"733ac18b" , x"1791d09e" , x"a3f5cf33" , x"0626a785" , x"f8ea2f52" , x"7dbbbb3b" , x"ee5f1c39" , x"473c81ec" , x"38dc8e87" , x"56fa534a" , x"a4e25bd6" , x"498fbe64" , x"bb15c0c4" , x"2bc05061" , x"f16ab5be" , x"66361ed5" , x"eaa685a2" , x"b299299c" , x"04c2f11c" , x"3424239d" , x"a37ab701" , x"aa945f75" , x"642af038" , x"716cc767" , x"dfcd18cb" , x"6eec7049" , x"19462537" , x"2cdc7df5" , x"d06eb82c" , x"3175b4f8" , x"542e066c" , x"9dcdc9df" , x"9fd63d0f" , x"44dde10c" , x"98bf07f3" , x"8f470d9f" , x"64aa7dd8" , x"f1dd5d0c" , x"d2f3df38" , x"b6e79cf4" , x"abb0da91" , x"ade156ca" , x"f5bdbf54" , x"f599f724" , x"e90d1dd6" , x"c67c4f25" , x"caa4e1ce" , x"9b93fe9a" , x"aa018231" , x"f2b0485f" , x"cef0cf82" , x"0f44ac6f" , x"363c6497" , x"44ca5518" , x"76cb48ab" , x"fc971022" , x"c416d981" , x"c5af5734" , x"20c24f3e" , x"79b0d1c1" , x"22a753f6" , x"ae4f6ee8" , x"57b8a79c" , x"6abc3c69" , x"87f84830" , x"6151755e" , x"5036a524" , x"3698e366" , x"124407bf" , x"62083958" , x"ddd13318" , x"07984e5c" , x"33daa03e" , x"78ea0892" , x"3dfbde8d" , x"5557e991" , x"9afd5eab" , x"f9d0f71b" , x"7cfdcf0d" , x"8e318c35" , x"c92bc43d" , x"d8a75ae4" , x"76215402" , x"6876d96f" , x"192e7620" , x"7646d294" , x"3c88e37a" , x"d388d64b" , x"b400df1a" , x"fdbf7e24" , x"7903b62c" , x"86216efa" , x"1339ea1f" , x"ece96e96" , x"bbd50e86" , x"bd30896f" , x"32202ba7" , x"91431883" , x"f034ed76" , x"f801d00c" , x"db7b159f" , x"d31264db" , x"dd8bc3e6" , x"f5a8f42b" , x"31df565d" , x"a576ef96" , x"67d7c390" , x"612bba58" , x"d3287e88" , x"7a00cc51" , x"e3dc7833" , x"e9719c50" , x"d1f82248" , x"03cd7655" , x"c5f0ad3b" , x"281d1693" , x"2ad59568" , x"78b8ac1c" , x"fc51a49d" , x"8b0180ea" , x"9ae141c8" , x"0f47e94c" , x"bfb13356" , x"a874ac89" , x"93989310" , x"e3bf23aa" , x"2b0a4b45" , x"1c10e1ff" , x"4eb87e74" , x"7011e61d" , x"c5143753" , x"47bd28ba" , x"f1bfb47d" , x"fc391a3a" , x"93dc3080" , x"9bd79c5d" , x"994082a6" , x"40f5b549" , x"08ce28e1" , x"21f309fb" , x"5640e6f8" , x"8b8570dd" , x"3f8b9a2f" , x"d3eaf55a" , x"e957baa9" , x"d6460b00" , x"04b833b8" , x"d556564f" , x"096df739" , x"3426b1ce" , x"bfdcca32" , x"8b5ef55f" , x"ad18ab53" , x"dffc3f11" , x"372e544c" , x"1ef9dc81" , x"a74b93fa" , x"db39cdc7" , x"862d1a93" , x"e657b896" , x"f9589fb3" , x"37c60221" , x"f1f8119f" , x"13b4e6aa" , x"e22bc29d" , x"79662a3f" , x"6c4bd791" , x"d5c45c3f" , x"44bcb2ab" , x"782a2c27" , x"61cbf5b5" , x"69ecd3ae" , x"2927e9e0" , x"80b3faa3" , x"4b601d99" , x"201cd555" , x"6e7b049b" , x"21dd7372" , x"d3a134e8" , x"ded77932" , x"ca097772" , x"9a5af162" , x"6e789398" , x"43ead05a" , x"e7c98ff8" , x"dd63b3b2" , x"76ba478e" , x"0ee042e1" , x"75483328" , x"752f5bc1" , x"710b102e" , x"b8e2bb3e" , x"921b1772" , x"56c8a5f6" , x"ebd0b5f2" , x"66b65829" , x"a008d4a0" , x"86e8252b" , x"0aa5d1de" , x"e4eca1ad" , x"e4528020" , x"c742a4ff" , x"1f96efcb" , x"11c21346" , x"06ec1c20" , x"475e6c45" , x"08771ed7" , x"611e61b0" , x"48864d63" , x"dd5b2e16" , x"a3b6a861" , x"6b8285c4" , x"a1e1585d" , x"3d689c31" , x"7d8ed6ae" , x"98ffe2ee" , x"526d7471" , x"7aba3f2f" , x"d83b45cf" , x"e6073590" , x"32470bfa" , x"ef491acb" , x"40df060a" , x"d1610810" , x"9861c3d1" , x"b57b0f0f" , x"81cae7ad" , x"be43b402" , x"5cd08a6a" , x"e653615e" , x"de66192c" , x"10b38e5a" , x"6178a0a2" , x"55fe4643" , x"3a5506f9" , x"011c1a78" , x"98a50431" , x"d3fe12c5" , x"6be77097" , x"81e748f0" , x"72cdf3b4" , x"5dbcd256" , x"424572fd" , x"3a050f6b" , x"fa0ed65f" , x"88eabb09" , x"eca8d78b" , x"4a1bae3a" , x"0ea4119a" , x"1180c141" , x"8433db40" , x"15c0a49b" , x"6a9d0d8d" , x"117eb20f" , x"254ae6fd" , x"68e9bbed" , x"69b37147" , x"1f95ec08" , x"cfa1ebe7" , x"71698915" , x"888ea907" , x"e620ea2e" , x"1ab12c11" , x"5a8815f6" , x"5a1373e7" , x"1ec3fe49" , x"29621237" , x"91b14281" , x"d0970ad9" , x"e0022502" , x"755b24e7" , x"593c35bc" , x"76ebdb84" , x"0abb55d6" , x"08c9f9cb" , x"2470602d" , x"bd8f46ff" , x"139b969f" , x"47379517" , x"bd932683" , x"56ed04c3" , x"74ded4b9" , x"5d1946d2" , x"ab12630b" , x"d6d63321" , x"b301ca66" , x"9492ff51" , x"9244775b" , x"ec6a8fe9" , x"a0f20bfb" , x"f74217d3" , x"e0b522f0" , x"bef68154" , x"a98fe22e" , x"a13585d7" , x"e01b1b5a" , x"0bcdd82a" , x"77af320e" , x"11de6b72" , x"242e991f" , x"9b9eba84" , x"1171428a" , x"0c5b8064" , x"b6d89730" , x"1918eea0" , x"4ed82c15" , x"f55dedbb" , x"abd166e8" , x"66097b97" , x"a7050d56" , x"3af0e484" , x"87f2d100" , x"8a2b03a4" , x"b711412a" , x"14784981" , x"813b44d3" , x"e475cd19" , x"7ced86a6" , x"29fdd1c2" , x"7f7254dd" , x"bfd69faf" , x"ef9c1815" , x"3b124590" , x"63a7f6f4" , x"0457e7d4" , x"1dfd39a2" , x"fd79bbdf" , x"3d8c65f5" , x"2bf4dce9" , x"af5629d3" , x"097a6b14" , x"d6d95320" , x"6dd88d4b" , x"f85b6606" , x"757ef1ce" , x"37155b0d" , x"90b0c1b3" , x"c2a5dc9f" , x"74c7bd1f" , x"9587c3a9" , x"6d200ca4" , x"6727d5a0" , x"3c521a05" , x"829200e6" , x"5279f281" , x"7ee28a17" , x"fb5fb9ed" , x"a6c0137d" , x"069665dd" , x"be6386aa" , x"07eb1695" , x"4d4cd284" , x"96858b66" , x"16f0cedf" , x"5831f51b" , x"d372794a" , x"7728528a" , x"63bbf96f" , x"321efdd6" , x"c67a60fb" , x"e9c20955" , x"2deb221a" , x"714325f6" , x"1bff18a9" , x"1982dc97" , x"e7b874f6" , x"9e713d20" , x"e0588a18" , x"ad4faef9" , x"fff267d7" , x"7897ec12" , x"dd3fcb96" , x"603d477a" , x"0970ce34" , x"41557e18" , x"8b704ee1" , x"d903293a" , x"ff63c625" , x"6382b696" , x"82d16e20" , x"73cf0994" , x"df9e7e63" , x"a269edff" , x"11fa08c4" , x"794c9a0c" , x"fccf56b4" , x"91acd7d9" , x"ec36f291" , x"1bdd659a" , x"9073674e" , x"a0bc46a2" , x"6e744c15" , x"8ff87008" , x"567cfb35" , x"f74385dc" , x"b88154b9" , x"00850a04" , x"037eee73" , x"21d1a897" , x"5fc268b5" , x"35a93439" , x"ec351929" , x"f0b1fff8" , x"8be61707" , x"c1b8f78a" , x"7950a649" , x"fcb6a957" , x"7f1d11c7" , x"bf8dab2c" , x"4f18ba87" , x"89f9f5bf" , x"f36a1702" , x"d83dcc75" , x"fb63e96a" , x"11ee4fe3" , x"8378df1a" , x"f12e5b9a" , x"fe1a5dd4" , x"4570e678" , x"74b22c46" , x"03a99d46" , x"6d1103f2" , x"118656f2" , x"36953e60" , x"2fafedbb" , x"3178cc58" , x"334d44f9" , x"d52f61cc" , x"e061bcbe" , x"ba04e39d" , x"96e8a7fb" , x"879d69f9" , x"742d52a3" , x"d43ea292" , x"ea6ceaa5" , x"830a33fc" , x"320d1a19" , x"8d4d5f16" , x"f26ca926" , x"3699d6a8" , x"e43b98cd" , x"967b698e" , x"efc34ccf" , x"248c2173" , x"bf88b022" , x"0d5e8574" , x"40b9e440" , x"aeed4465" , x"eab20792" , x"9bca8dd6" , x"8b99b348" , x"383b5f1b" , x"820f2538" , x"6801f659" , x"c9a3edcc" , x"a141a5aa" , x"31f6a2a8" , x"8e28a3f6" , x"bb527595" , x"20a9056f" , x"d8de9ad5" , x"2b5094ef" , x"a7fd2df2" , x"00417f61" , x"a1030b09" , x"6b0cb210" , x"d1a64580" , x"7d0d65a9" , x"fab5a1d9" , x"28ed2a08" , x"e7e9e8f9" , x"aab5eed6" , x"c719039f" , x"04966dfe" , x"380f2429" , x"1ea30b55" , x"7319288a" , x"f3be7bf6" , x"ba99596f" , x"f9d190c8" , x"d69a9fdc" , x"07ea03f5" , x"2469f1bc" , x"7e6f0a53" , x"f812d39c" , x"dcdb5b64" , x"ef22658f" , x"3e2d21e0" , x"39a7747d" , x"d592bab1" , x"e99b410d" , x"d0478334" , x"5d78c18d" , x"a10461bf" , x"008c29a5" , x"0092aeb4" , x"ecf74315" , x"6135968b" , x"75156b58" , x"e78721b7" , x"c6024691" , x"ae2b86da" , x"b9db1145" , x"60fa8d71" , x"eb7f73a2" , x"a1c7c8b8" , x"782846d5" , x"3e46e95d" , x"98ff6dc7" , x"92482082" , x"385d79ec" , x"fb5293a5" , x"874b9b9a" , x"d984c2de" , x"19966c24" , x"488fcc4d" , x"9e34f986" , x"aeb58bae" , x"2dbeee95" , x"5bae0c8a" , x"e3b44961" , x"fca73b8b" , x"c443b620" , x"15802020" , x"ccae1c1e" , x"40140bfb" , x"5f5bbe18" , x"cfb46974" , x"53fc66af" , x"159cc0b7" , x"31772b28" , x"88004289" , x"01221751" , x"ccf5a0a2" , x"3eeeaab5" , x"bd23850d" , x"ec9af5c2" , x"2444067f" , x"5b9fa606" , x"7019d687" , x"667752ae" , x"59b2873e" , x"8568c1df" , x"7a7ecfcd" , x"ed7496e3" , x"966011ba" , x"c8bccc3c" , x"255385a1" , x"244e9e43" , x"e7c3bf31" , x"31757b14" , x"a3e3c520" , x"7d64c105" , x"29b66876" , x"147ed6ab" , x"90df843e" , x"c67f48ae" , x"ee7e6537" , x"45f179b3" , x"c8795d76" , x"9ee4532b" , x"af893136" , x"a4e6aa2f" , x"775a25b0" , x"2e1f809d" , x"42a434f9" , x"5b8ed623" , x"91bb8f10" , x"8b6fad99" , x"3faf6f38" , x"2a77df2a" , x"51bdbfc4" , x"2924df1e" , x"e92a55de" , x"43f6e6cd" , x"e29dc7cc" , x"aead9d57" , x"cb6a3672" , x"3451866c" , x"ed01df09" , x"e0c84d6e" , x"2dc87472" , x"de67b90c" , x"847d93b0" , x"1014498f" , x"a0836bb6" , x"032b3f31" , x"e9c65178" , x"b76e7a57" , x"a9f9d2da" , x"7e8f2b29" , x"63a22415" , x"74bac1f3" , x"bd712311" , x"47cba27a" , x"d15084b1" , x"3425fc2a" , x"99b0325c" , x"2822a7db" , x"15c25e0a" , x"e25c636f" , x"ec1fa77c" , x"4f15f1e7" , x"0db89611" , x"ff5f9215" , x"86eb1b6f" , x"bf66e167" , x"1e6d2b0c" , x"c0d58514" , x"61510d1d" , x"771c2fc8" , x"d015cae9" , x"d365db17" , x"3e7d11f4" , x"33bd9d81" , x"e26985ff" , x"e52fa38b" , x"b670052f" , x"a8b7da86" , x"60ce561e" , x"34c531c4" , x"3fb93217" , x"a47c0ecd" , x"40bb05e9" , x"33ca5463" , x"c46a139e" , x"1478285d" , x"0cc3bf9e" , x"ecc22b37" , x"af6f1258" , x"919fa401" , x"9eca8c0e" , x"4880b447" , x"bf26b944" , x"9121dd8b" , x"fa2d6d04" , x"cbceb2ba" , x"624827e8" , x"6af566c9" , x"429cd598" , x"c16329f7" , x"e0a1d7ef" , x"8355ed5b" , x"ce5c4e69" , x"74ebe4c9" , x"760c07f7" , x"a9333bb8" , x"174943e2" , x"16968123" , x"9073ebf5" , x"b59b1542" , x"2ff8533c" , x"a5c93c66" , x"881ccf17" , x"3855518d" , x"5ae376aa" , x"d00e2dc2" , x"5095a6c3" , x"d1f5fac4" , x"ba0bba9a" , x"ca9c6947" , x"8409b0b7" , x"2ec8b16a" , x"ca67b434" , x"da444dc4" , x"3459a03f" , x"a9b0d18a" , x"ad985c2f" , x"12b48e29" , x"0d6fb15e" , x"49251eef" , x"cd19a1d7" , x"3672ad06" , x"adb6ac9c" , x"fe8fbf6b" , x"f22da470" , x"46e04540" , x"17705abe" , x"eaa39dfe" , x"e88f6ada" , x"2084b7de" , x"828c4849" , x"051d7762" , x"9d6a51e0" , x"73c342f1" , x"50ea0ac2" , x"7819e4e9" , x"13d63839" , x"b7aa45d4" , x"d9c1d7e0" , x"58072e10" , x"24ffb728" , x"15e31c8f" , x"5ed82820" , x"58a7279e" , x"9f550b8c" , x"132807ad" , x"ff5f8fa4" , x"e80ae452" , x"8470aa4f" , x"288aaec7" , x"fd92249e" , x"db2274e0" , x"39fe2981" , x"e0c10d46" , x"65e3aaf4" , x"da81706c" , x"b2525352" , x"e6f5e839" , x"108c4be0" , x"debb5b72" , x"bf66bfcc" , x"e65350ea" , x"6b9f5cdf" , x"baf42ea6" , x"cfb27f99" , x"d4c77932" , x"612dcfd9" , x"fe302631" , x"51ae6da6" , x"e84bf945" , x"fc6dd7a9" , x"de36ba52" , x"b7dab43e" , x"63e64eb9" , x"69c66267" , x"a2792428" , x"193fd4cb" , x"5ad71d09" , x"bc0c110b" , x"dc8b77e4" , x"a326815c" , x"54d388d5" , x"12e74d04" , x"ed40dad3" , x"1ed99f9c" , x"4cc785f2" , x"fb49e383" , x"f9633863" , x"7f2e3f2d" , x"a9b48b4b" , x"05bce6aa" , x"c66f3660" , x"0dc7e78b" , x"32895caf" , x"24104e23" , x"0c817f0b" , x"e4babb90" , x"25ebf13a" , x"773ffbfc" , x"ded47d48" , x"8f944ebd" , x"2032cabe" , x"7e94b0e0" , x"8a7d91ec" , x"115a63c6" , x"41850a2b" , x"e5cc29fd" , x"76e65d2d" , x"49df6a95" , x"233dc1a3" , x"44e04096" , x"33acb2e4" , x"981d1c1e" , x"3793a694" , x"79d33533" , x"6964d808" , x"5e49a1df" , x"ba3fa4d5" , x"a7d620f2" , x"049e7031" , x"f02de6cd" , x"e02f96c3" , x"9ed42f4d" , x"d474b22c" , x"48683549" , x"7bd97089" , x"3486c222" , x"766fa555" , x"706b1752" , x"b808d1dd" , x"06f9decf" , x"920424c9" , x"e04d9dd9" , x"e1bcc066" , x"9c2f0174" , x"2a55f057" , x"341ea15e" , x"b864e237" , x"851944d1" , x"f8eb637b" , x"0dc76de0" , x"8bb7e3a2" , x"dcb850cd" , x"1d5a9d82" , x"71642a8f" , x"87ba78f3" , x"8c4a540c" , x"0552459f" , x"911dca9b" , x"ef585dc9" , x"ae2e5dbb" , x"dd056ea9" , x"5f12aa89" , x"fac22ce2" , x"1406cbfa" , x"9c7c8b06" , x"74d366a4" , x"4ca996df" , x"0c3f7dc3" , x"2809ec41" , x"bcfe6908" , x"26631c82" , x"09ba77ea" , x"bdc99a31" , x"f4495b2d" , x"2c236fc7" , x"be0c1d0a" , x"0fcfab85" , x"effcb1f3" , x"00b6df21" , x"836bd260" , x"dbee3a9c" , x"3dabefd3" , x"cbe8059d" , x"428d15ae" , x"1179cc76" , x"c24c2166" , x"8bc93189" , x"fe4bb61c" , x"e35719d8" , x"5b51117e" , x"51c4f204" , x"c0bb4a9f" , x"f098c36a" , x"1c2c2378" , x"40953419" , x"98d7f4d5" , x"3b69d357" , x"6e3b7cb5" , x"79885089" , x"bb10560a" , x"17f41ad0" , x"42dc7102" , x"38c8d24d" , x"184550e4" , x"9e7ce796" , x"737257c4" , x"f190a4f5" , x"a3dbec42" , x"84d348f3" , x"21cd4bcd" , x"13366fe5" , x"73ec2ba2" , x"b7ea9ca6" , x"a6f68d8d" , x"5f929fb0" , x"d3b629bd" , x"1f1b8ca5" , x"4ede20dc" , x"b28a70fb" , x"67014cb4" , x"676cfe50" , x"e25cfbd4" , x"4425f5e6" , x"b3592ddd" , x"1f79efdd" , x"3deb57bb" , x"ebbd2038" , x"c2845676" , x"f7ceb353" , x"4a7a1bfd" , x"767bd873" , x"4706395a" , x"8476ba51" , x"019047f7" , x"71ff49f7" , x"5fed11c8" , x"055609f5" , x"6fdad3b7" , x"1e5a9379" , x"4de68126" , x"1f2edcbe" , x"4a75d287" , x"bd5b48aa" , x"3e158c6b" , x"fb42fe62" , x"efca7f2a" , x"fdf60e74" , x"dc356d6b" , x"c5861dfa" , x"65b0c047" , x"9d051120" , x"7abb35d0" , x"f26206e8" , x"90a3957a" , x"f1ae79d2" , x"7d57b24f" , x"0cb81c2e" , x"45126010" , x"5350b310" , x"fd5f9c3b" , x"2d909be5" , x"2f055ecc" , x"a443a67c" , x"dc9588f0" , x"ef6acb4d" , x"085a9ba3" , x"afda4c86" , x"54fb3361" , x"2e282455" , x"bfade21a" , x"9eedac29" , x"a4f5335a" , x"043c70a4" , x"2b532dde" , x"d6a5015f" , x"f3c3b6ac" , x"357f77e6" , x"8b13c21f" , x"af330fa1" , x"405ca22b" , x"8ee742ea" , x"941d5091" , x"e98a1cfa" , x"ea5cacb7" , x"28d028ed" , x"e545d047" , x"f19c708c" , x"7b858dbf" , x"ee01bf70" , x"71576820" , x"e9041e46" , x"4fcf2c23" , x"622e2233" , x"0e290b19" , x"cd6ff36f" , x"c0f87f6d" , x"36462a8a" , x"21c74f44" , x"f2e6f30f" , x"5b1db642" , x"2b16d639" , x"6557ccb2" , x"5f087860" , x"e2b184f2" , x"3fdaa475" , x"056ff465" , x"f5b45ff1" , x"d815ac93" , x"6173915f" , x"49beff6c" , x"513bb992" , x"40167896" , x"ea3e7ec0" , x"7d0672a3" , x"03b796ed" , x"baa21c66" , x"0813e5bc" , x"33dea619" , x"1555623a" , x"375de08a" , x"ea05b486" , x"f9f10f00" , x"577816fb" , x"97de4d04" , x"3aa72eee" , x"4ded6492" , x"a59318ff" , x"f7bb6041" , x"5c8cffff" , x"e55e4766" , x"06cfde8d" , x"30a58275" , x"c1d652a9" , x"0075ebb7" , x"29ba2465" , x"b6362672" , x"2f55f08f" , x"de2357d3" , x"21d917b3" , x"1e496d40" , x"dce6015b" , x"09fd68e7" , x"46b3cd92" , x"992346c6" , x"1aefe4f2" , x"9ab44a33" , x"b9bdc804" , x"8434ea15" , x"cbc78526" , x"01ec015e" , x"b877d4c6" , x"b05defd4" , x"cddfba5f" , x"f22e642b" , x"6d5c6c64" , x"dfa015d1" , x"83053410" , x"1cffaf83" , x"17faacb8" , x"5ac50e72" , x"64b0697c" , x"3def9277" , x"b9eaa4bb" , x"8f7200e0" , x"c4ffc5e3" , x"9cdbaf06" , x"42653aeb" , x"4d01d318" , x"b5d18970" , x"cc5303eb" , x"8055260a" , x"cbaf2b66" , x"7104fbdc" , x"c7f5a9a8" , x"49f2fd77" , x"59e1963f" , x"e72e3b1f" , x"0de66e64" , x"7a13f278" , x"b56daa77" , x"83998d9b" , x"fe308ef8" , x"7559f25a" , x"29980f0e" , x"b213a527" , x"1d12aee0" , x"f42ee73c" , x"e9b23439" , x"9c09c806" , x"7b4ddf26" , x"94b8cf35" , x"da0ff473" , x"934febe6" , x"cf5682d4" , x"874ad847" , x"2fcf7935" , x"b6d6b029" , x"3f487d60" , x"226358b5" , x"0ddf51ef" , x"2bd82cfc" , x"9be4e5e0" , x"1ff394ae" , x"c6f8b441" , x"c79f7349" , x"82d51891" , x"e7317fbc" , x"071aa134" , x"d2c57f8b" , x"fd89e3d6" , x"5627e643" , x"803d9947" , x"6e427ea3" , x"54fdc990" , x"66d19eb4" , x"2c839afb" , x"fb197d73" , x"a029b4fb" , x"78813eba" , x"933c0954" , x"8d8c7e5e" , x"c040940d" , x"127c7477" , x"274d0201" , x"82e492e3" , x"5b5667de" , x"e84f290c" , x"24d9f5ac" , x"5a526007" , x"d9c16c59" , x"e80b7065" , x"567ea188" , x"e7756a46" , x"46734710" , x"05f507a5" , x"0189ef77" , x"27a42563" , x"cd4a1a50" , x"7bdd7490" , x"7f562620" , x"ddb164be" , x"89b01180" , x"2effa07b" , x"def41f98" , x"57673003" , x"b90c46b7" , x"7c5edf83" , x"ab07adfe" , x"dbb0705a" , x"2dc7a86d" , x"fc7b82cc" , x"8ced4379" , x"ce4a60e7" , x"f5ba5f9c" , x"39ae9f58" , x"9894e059" , x"a71b6ed2" , x"cefe7d74" , x"74c2a72e" , x"fc0a4fea" , x"cff05b78" , x"e2cbf1ce" , x"8bc10404" , x"36be0595" , x"b85d1cb2" , x"08dd8414" , x"265d3961" , x"737cd949" , x"54317ae3" , x"03880a5d" , x"11cc407e" , x"79451b96" , x"7a50e89e" , x"f381a709" , x"65d81a6f" , x"3fbb5636" , x"3a6fa4f8" , x"62ec9ace" , x"567ac803" , x"6e726aeb" , x"9138d9fe" , x"d4b4fa15" , x"357bf7a5" , x"d31c0dd7" , x"88966816" , x"73f7b78e" , x"87bbb7ef" , x"616c643c" , x"60af0f40" , x"ed05b898" , x"3f2a635e" , x"bda7ed8a" , x"7ad278b0" , x"bcd58561" , x"36645c59" , x"f2691625" , x"fe86d1ae" , x"8295e4f2" , x"84401eff" , x"cab89831" , x"0c1e117d" , x"73c1a489" , x"24f7fcf9" , x"d9651631" , x"25d3ab0f" , x"63f3464b" , x"df21f58b" , x"bd063e3c" , x"c86ebbc8" , x"f9f7e084" , x"b3097943" , x"85f6ed5e" , x"a87df30d" , x"6e0eeded" , x"0725cbd1" , x"35084ffc" , x"2e7d9b88" , x"52ca6ec7" , x"62ae794c" , x"1c61fd90" , x"cfa80b30" , x"600dc427" , x"00cd5349" , x"5474964d" , x"899b8c33" , x"57943445" , x"f2f25be1" , x"d12eb37e" , x"ba792043" , x"881c8744" , x"e34f82e4" , x"8568413d" , x"5c8fb5b8" , x"c639293c" , x"e8956037" , x"1ec98a6b" , x"db692b9d" , x"a01d804a" , x"5e1cad09" , x"58bdf7c7" , x"fd20bd1e" , x"55a99da3" , x"b651a730" , x"931a123c" , x"9bb089b1" , x"dd2b0461" , x"510bff37" , x"32d5079b" , x"6954765f" , x"ac25bf0d" , x"89f5ee27" , x"e6de6ba2" , x"a6ee160e" , x"32fbf707" , x"6e8914c7" , x"4c5c599a" , x"e37ac19a" , x"7f1bf3cf" , x"94a88122" , x"e3d0c394" , x"1d42fbd7" , x"805cb4fb" , x"09c8760d" , x"46e928ea" , x"a8cb4fb7" , x"88b17bac" , x"96725e4c" , x"930204d6" , x"6a03f095" , x"69ad8c93" , x"e84b5a87" , x"03c78d34" , x"4755ab3c" , x"b3e864f6" , x"3c08a635" , x"81ba2e7d" , x"57d280aa" , x"619aa7a5" , x"7e89da79" , x"109f5a6f" , x"16192c1b" , x"5bcbe574" , x"a051f8d0" , x"3bf7e3bd" , x"8dc969f8" , x"3418d768" , x"9e17b76c" , x"d053dbd2" , x"bebe2128" , x"64b8213f" , x"44cac8ea" , x"0db71a3f" , x"b5d26332" , x"6003615c" , x"b7f28f18" , x"c66604aa" , x"b4cb6f76" , x"2a50f1eb" , x"1df9066a" , x"e9872d69" , x"cc86706b" , x"51b7785c" , x"cc84a493" , x"546c70a6" , x"d152826a" , x"3448c9e6" , x"9de19016" , x"c4682f4f" , x"ce15a06f" , x"11e9c2b5" , x"12cdddda" , x"f3356cdd" , x"067745ae" , x"28806fad" , x"e0a87c79" , x"49548439" , x"6222317a" , x"afe7b186" , x"9f65a614" , x"24226507" , x"a2e243af" , x"83181c44" , x"c45b30ba" , x"b8a8e1b8" , x"539ef063" , x"edc8cb66" , x"c449a6f9" , x"bb6b2863" , x"68c3a378" , x"bff60a25" , x"b053165f" , x"684618e4" , x"b2dcdd3b" , x"3d4f53e0" , x"41b5575e" , x"855674ea" , x"64b3a458" , x"38157426" , x"87b1ad1e" , x"d7a6bbc6" , x"8e543136" , x"a9b5f89d" , x"de8a23e3" , x"d0f4cbad" , x"7d0c9ced" , x"cb3b8ff7" , x"cbbd74e9" , x"7817474b" , x"9d1b1df6" , x"4f3d0765" , x"7c4bec82" , x"b0053188" , x"6bd6a6f6" , x"fca258fa" , x"4b8ef1c1" , x"c51a62f8" , x"870e7e1e" , x"d45f690c" , x"7094df03" , x"b4c1f880" , x"fe80dd10" , x"9867f7b7" , x"81adc38b" , x"c0bc5bbe" , x"de13095b" , x"7f292fa4" , x"a502f680" , x"dd795572" , x"3d77c69e" , x"116a4348" , x"8c109fe9" , x"f7f2a06e" , x"8f1b64b0" , x"194817fd" , x"d1831c5d" , x"8c06b0ac" , x"cfe4e7c0" , x"67290922" , x"a2b6ac16" , x"1b66fbcd" , x"766b9b48" , x"b962f459" , x"18abb12b" , x"9d1a4946" , x"74fc3d8b" , x"c8709a70" , x"e562f176" , x"910e0be8" , x"369e5ff1" , x"cfb29cda" , x"2a1da0d5" , x"93a79522" , x"86dbcadf" , x"f1abe5a3" , x"90274e83" , x"df177ce7" , x"7dde0eb2" , x"81f237f9" , x"14005ac7" , x"c9f050a1" , x"0072231a" , x"79188934" , x"e55c6d1f" , x"d42c590e" , x"ef045019" , x"528e2757" , x"124e4c6f" , x"f9e4bd5b" , x"273ddbfc" , x"4738d6a2" , x"ba87ddfc" , x"12a50a30" , x"267c662f" , x"c05030a5" , x"99a0b391" , x"d4c8c711" , x"30034b4c" , x"ec1e597b" , x"55b2982e" , x"53b7dd34" , x"a82c7ce5" , x"cdd77ba6" , x"93ae2cf6" , x"89cac609" , x"d4b23f86" , x"769a7e46" , x"1066319c" , x"d21cb028" , x"ecd63ada" , x"f3b02508" , x"87890b1a" , x"13869ea4" , x"edb8d23c" , x"b56b7789" , x"22773f02" , x"3c2423a3" , x"89f6ab4c" , x"661e04ea" , x"7761f83c" , x"44a3cd70" , x"6694be73" , x"d51f97a0" , x"e2193b6f" , x"fed0d164" , x"55dad64f" , x"a6561483" , x"abcce151" , x"b43640bf" , x"9a1810c4" , x"eeab6c34" , x"09db312c" , x"b009ff5c" , x"a7c1d4b3" , x"917fa466" , x"a9ed407b" , x"617f395a" , x"187cc435" , x"a273cd1d" , x"afc94cd4" , x"5cfc8d0a" , x"448edc35" , x"6859bf62" , x"ca0cf9eb" , x"5e631afb" , x"366b07b2" , x"77e8fb30" , x"6ae880e4" , x"80dfbac9" , x"4a10f821" , x"e918df75" , x"f9ebff8b" , x"34d8a9c2" , x"c57eb17c" , x"56aebaf0" , x"fcf95f21" , x"92f9e597" , x"91e29e97" , x"7ca79abd" , x"b5b1d43f" , x"4320c891" , x"7f72260b" , x"94603cb2" , x"c2df4d22" , x"e0da1586" , x"3229cf65" , x"0f9a6f0e" , x"5e9a4232" , x"70dd47b5" , x"fd0ca72e" , x"1591eea1" , x"815d9761" , x"90305721" , x"110b5319" , x"8a104210" , x"c5e99fe7" , x"c49f7153" , x"58cc1e14" , x"3babcdd8" , x"c0e1a4f9" , x"965d56c5" , x"973529c7" , x"757f4fa7" , x"9dc3fcbe" , x"dc6948fe" , x"b4db6ee9" , x"a92c8de3" , x"2d5f6390" , x"5a97d32c" , x"a95f5922" , x"58e13381" , x"18969b6b" , x"40f3ab70" , x"3ec03e8b" , x"f3d8e265" , x"872faa5c" , x"4c56e67d" , x"576dd67a" , x"288d4ce5" , x"dc5cff35" , x"5c7df6df" , x"164576d9" , x"bddb676e" , x"dd8d0fb7" , x"b4b5dcf6" , x"8a947109" , x"b36dab79" , x"0407757a" , x"01980368" , x"0a980f1b" , x"5fd51d06" , x"170caf24" , x"e6c86aaf" , x"d2cb3c19" , x"517f0bec" , x"8b8a535b" , x"98da6d3b" , x"61a955f4" , x"4c3c4e05" , x"ccffecce" , x"2000f142" , x"39370ab5" , x"636b46e5" , x"80c941e4" , x"d153fbea" , x"35a98674" , x"fb2e54b1" , x"cad6beff" , x"dcab5db5" , x"405790b7" , x"15754913" , x"5a97ff9c" , x"56744b00" , x"0fb85ac2" , x"3c72f608" , x"3999cd1b" , x"515bb1b8" , x"1d4a4583" , x"fc04cf8e" , x"50e4b915" , x"8c5a2b83" , x"ff97e27f" , x"bfceee3e" , x"bb500784" , x"d783986e" , x"25c44296" , x"2ab948a2" , x"4c62f009" , x"e73167b6" , x"47f4d561" , x"1ae96a3f" , x"9822b862" , x"bebe6bc5" , x"8d819a0c" , x"bab81e91" , x"5d12537c" , x"b7ac1663" , x"e780a163" , x"22289586" , x"b540a2d4" , x"721f3a4d" , x"aeb621d5" , x"823fe14f" , x"35830321" , x"87ce362e" , x"8f4b6146" , x"dc166a95" , x"501b9e55" , x"ad7f612d" , x"b9cdfe47" , x"ce4b6a83" , x"3b1cc3b9" , x"87ff8846" , x"f4766282" , x"f4b596ed" , x"a9cf29e5" , x"1111bd92" , x"039c41b9" , x"8aa0ecf7" , x"50bc5993" , x"481ae46c" , x"5f1de2c5" , x"7b1c48c5" , x"8a9a305c" , x"af533b84" , x"b8dd34dd" , x"35506bea" , x"c7ff5ab2" , x"9bb0705b" , x"25b76267" , x"5380481d" , x"c8bdc000" , x"e17f33da" , x"375622c3" , x"2226262d" , x"eec82ab8" , x"1a376587" , x"e35fc221" , x"f588af63" , x"a0021feb" , x"272495ed" , x"00c51722" , x"270cbc5b" , x"ad98b146" , x"27d24b4f" , x"f4174cfa" , x"16ee052d" , x"c2584cad" , x"74552b12" , x"2dcdfe57" , x"ab3cbf80" , x"28718ed2" , x"d4d02fe4" , x"08b32799" , x"ca4cd981" , x"a98e4c81" , x"b6743900" , x"1b598fcb" , x"78fc2662" , x"629aeb91" , x"b566087c" , x"e6fb80b1" , x"f54362de" , x"d4d691b1" , x"817a81d1" , x"d97c44d4" , x"4e17f615" , x"0ea6e2c9" , x"ca3110c8" , x"a38e56cd" , x"3c83db30" , x"2e7bddbb" , x"3bfb453a" , x"f2249978" , x"76f68a27" , x"7bf69d35" , x"9e902225" , x"365f5c6f" , x"9d863a5c" , x"0fe514ca" , x"1f6447a6" , x"772116bf" , x"1fb0eed1" , x"1cf97f34" , x"48d24dfd" , x"8559783e" , x"bc58fc24" , x"bf4cb705" , x"694b7ce0" , x"1722b4e0" , x"d438285b" , x"316b164f" , x"ef63a383" , x"13b15028" , x"66293b85" , x"2dd702af" , x"0d5db981" , x"d11e6789" , x"9239408d" , x"e85a015d" , x"bf674cb2" , x"6e08b7ac" , x"51fb7b5d" , x"c67f8c3b" , x"7e30f18e" , x"4d27794e" , x"38be3c29" , x"1c5714f7" , x"f0743e65" , x"b59a400a" , x"7b785c0f" , x"23d7f1ba" , x"8a3d2eec" , x"e8bb8c12" , x"389732b4" , x"ae34a9bc" , x"188fda08" , x"284ac302" , x"0f670024" , x"80597501" , x"d1cb5572" , x"4545388d" , x"c57f9a3e" , x"42f98e48" , x"32191d97" , x"6592994a" , x"e526769c" , x"fee4bd54" , x"af2e4b44" , x"e5721d24" , x"a8271747" , x"5b9c093d" , x"fd899f46" , x"b7b629f6" , x"08a00671" , x"ecc96881" , x"6c9bdcd8" , x"0d8ad067" , x"7d6f91e7" , x"5236ef43" , x"95608c84" , x"4dd06639" , x"15512a9f" , x"54dcd80f" , x"a8ffe4d4" , x"9075e2e3" , x"0d63dff9" , x"e4f38018" , x"8e8c7237" , x"2c16ccef" , x"b6474967" , x"37afcbbf" , x"7ce7b5fb" , x"96e7414b" , x"9e1b136d" , x"813cbc2b" , x"36ba2082" , x"61c4da5f" , x"a549e2d5" , x"af760cbc" , x"6171c5fd" , x"8455f8f7" , x"1a8cecb0" , x"c63943a2" , x"60a49856" , x"5798246e" , x"434ad884" , x"5d32d2ac" , x"3dc4e4dd" , x"bab83ef3" , x"9f77f346" , x"c200cedf" , x"85de981b" , x"2518def9" , x"69c9f2fa" , x"75526191" , x"37c13809" , x"2f4d8b66" , x"dbca2b79" , x"db2bf71d" , x"dc6b0974" , x"8c1068b6" , x"48b03a2f" , x"05d60bc2" , x"9d8a62dc" , x"034ae867" , x"c78c9fb9" , x"eff62aa4" , x"f470df89" , x"b9c27935" , x"eb6b1e46" , x"5eb2a304" , x"6283482c" , x"6dff30c2" , x"29a2f902" , x"231a17b1" , x"cbf7e6a5" , x"57d3810a" , x"1d231f61" , x"42033023" , x"28a8b58c" , x"84f7ef8c" , x"5b178d37" , x"52696449" , x"d906b49b" , x"67de50c6" , x"9531261a" , x"2e54ded4" , x"960fbd42" , x"6ed031a8" , x"ed03b7eb" , x"5f78bd1b" , x"93385457" , x"838dbf39" , x"028de0f4" , x"486d4a0b" , x"cf33599c" , x"65b43515" , x"9bdadd50" , x"cfcdaf75" , x"7adb9f62" , x"d0f37879" , x"44b87e98" , x"26587765" , x"42129adf" , x"43d3732d" , x"7b2370f1" , x"0f08a8c9" , x"3a330d2d" , x"75a5a099" , x"0c713354" , x"0bacc78c" , x"2b536e7c" , x"d498fd1a" , x"42298993" , x"3c7cbcdc" , x"32aa3bd5" , x"460688ba" , x"9b0eb35d" , x"f0a40d0f" , x"d2de3def" , x"d4059c63" , x"cf847640" , x"929518b5" , x"cd5f67b4" , x"9be9dd90" , x"b546eb0f" , x"8c37881a" , x"dc002fff" , x"191af2df" , x"c7f527af" , x"61d2a893" , x"342c07c8" , x"5235810f" , x"fe4bbe5f" , x"213ec560" , x"17f7c6fe" , x"767623d7" , x"a68eefc9" , x"c209e291" , x"3715cf18");
end package;

package body utils is
   -- Taken from https://stackoverflow.com/questions/12750007/vhdl-use-the-length-of-an-integer-generic-to-determine-number-of-select-lines 
   function f_log2 (x : positive) return natural is 
   variable i : natural;
   begin
      i := 0;  
      while (2**i <= x) and i < 31 loop
         i := i + 1;
      end loop;
      return i;
   end function; 
   
   function muxSelectFromRand(rand: std_logic_vector(31 downto 0); numEntries: integer) return integer is
   constant increments : unsigned(31 downto 0) := x"3FFFFFFF";
   variable i : integer;
   begin
        i := 0;
        while(increments * i > unsigned(rand)) loop
            i := i + 1;
        end loop;
        return i;
   end function;
   
	function bitAdderTree(v: std_logic_vector) return natural is
		constant size: natural := v'length;
		constant vv: std_logic_vector(size - 1 downto 0) := v;
		variable h: natural;
	begin
		h := 0;
		if size = 1 and vv(0) = '1' then
			h := 1;
		elsif size > 1 then
			h := bitAdderTree(vv(size - 1 downto size / 2)) + bitAdderTree(vv(size / 2 - 1 downto 0));
		end if;
		return h;
	end function bitAdderTree;
    
   -- code de https://vhdlwhiz.com/random-numbers/
   impure function rand_slv(len : integer; seed: integer) return unsigned is
      variable r : real;
      variable slv : std_logic_vector(len - 1 downto 0);
      variable seed1, seed2 : integer := seed;
    begin
      for i in slv'range loop
        uniform(seed1, seed2, r);
        slv(i) := '1' when r > 0.5 else '0';
      end loop;
      return unsigned(slv);
    end function;
end package body;